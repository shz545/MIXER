`timescale 1 ns / 1 ps

module dense0_stage0 (
    input [511:0] inp,
    output [1394:0] out
);

    // verilator lint_off UNUSEDSIGNAL
    // Explicit quantization operation will drop bits if exists

    wire [7:0] v0; assign v0[7:0] = inp[7:0]; // 0.0
    wire [7:0] v1; assign v1[7:0] = inp[15:8]; // 0.0
    wire [7:0] v2; assign v2[7:0] = inp[23:16]; // 0.0
    wire [7:0] v3; assign v3[7:0] = inp[31:24]; // 0.0
    wire [7:0] v4; assign v4[7:0] = inp[39:32]; // 0.0
    wire [7:0] v5; assign v5[7:0] = inp[47:40]; // 0.0
    wire [7:0] v6; assign v6[7:0] = inp[55:48]; // 0.0
    wire [7:0] v7; assign v7[7:0] = inp[63:56]; // 0.0
    wire [7:0] v8; assign v8[7:0] = inp[71:64]; // 0.0
    wire [7:0] v9; assign v9[7:0] = inp[79:72]; // 0.0
    wire [7:0] v10; assign v10[7:0] = inp[87:80]; // 0.0
    wire [7:0] v11; assign v11[7:0] = inp[95:88]; // 0.0
    wire [7:0] v12; assign v12[7:0] = inp[103:96]; // 0.0
    wire [7:0] v13; assign v13[7:0] = inp[111:104]; // 0.0
    wire [7:0] v14; assign v14[7:0] = inp[119:112]; // 0.0
    wire [7:0] v15; assign v15[7:0] = inp[127:120]; // 0.0
    wire [7:0] v16; assign v16[7:0] = inp[135:128]; // 0.0
    wire [7:0] v17; assign v17[7:0] = inp[143:136]; // 0.0
    wire [7:0] v18; assign v18[7:0] = inp[151:144]; // 0.0
    wire [7:0] v19; assign v19[7:0] = inp[159:152]; // 0.0
    wire [7:0] v20; assign v20[7:0] = inp[167:160]; // 0.0
    wire [7:0] v21; assign v21[7:0] = inp[175:168]; // 0.0
    wire [7:0] v22; assign v22[7:0] = inp[183:176]; // 0.0
    wire [7:0] v23; assign v23[7:0] = inp[191:184]; // 0.0
    wire [7:0] v24; assign v24[7:0] = inp[199:192]; // 0.0
    wire [7:0] v25; assign v25[7:0] = inp[207:200]; // 0.0
    wire [7:0] v26; assign v26[7:0] = inp[215:208]; // 0.0
    wire [7:0] v27; assign v27[7:0] = inp[223:216]; // 0.0
    wire [7:0] v28; assign v28[7:0] = inp[231:224]; // 0.0
    wire [7:0] v29; assign v29[7:0] = inp[239:232]; // 0.0
    wire [7:0] v30; assign v30[7:0] = inp[247:240]; // 0.0
    wire [7:0] v31; assign v31[7:0] = inp[255:248]; // 0.0
    wire [7:0] v32; assign v32[7:0] = inp[263:256]; // 0.0
    wire [7:0] v33; assign v33[7:0] = inp[271:264]; // 0.0
    wire [7:0] v34; assign v34[7:0] = inp[279:272]; // 0.0
    wire [7:0] v35; assign v35[7:0] = inp[287:280]; // 0.0
    wire [7:0] v36; assign v36[7:0] = inp[295:288]; // 0.0
    wire [7:0] v37; assign v37[7:0] = inp[303:296]; // 0.0
    wire [7:0] v38; assign v38[7:0] = inp[311:304]; // 0.0
    wire [7:0] v39; assign v39[7:0] = inp[319:312]; // 0.0
    wire [7:0] v40; assign v40[7:0] = inp[327:320]; // 0.0
    wire [7:0] v41; assign v41[7:0] = inp[335:328]; // 0.0
    wire [7:0] v42; assign v42[7:0] = inp[343:336]; // 0.0
    wire [7:0] v43; assign v43[7:0] = inp[351:344]; // 0.0
    wire [7:0] v44; assign v44[7:0] = inp[359:352]; // 0.0
    wire [7:0] v45; assign v45[7:0] = inp[367:360]; // 0.0
    wire [7:0] v46; assign v46[7:0] = inp[375:368]; // 0.0
    wire [7:0] v47; assign v47[7:0] = inp[383:376]; // 0.0
    wire [7:0] v48; assign v48[7:0] = inp[391:384]; // 0.0
    wire [7:0] v49; assign v49[7:0] = inp[399:392]; // 0.0
    wire [7:0] v50; assign v50[7:0] = inp[407:400]; // 0.0
    wire [7:0] v51; assign v51[7:0] = inp[415:408]; // 0.0
    wire [7:0] v52; assign v52[7:0] = inp[423:416]; // 0.0
    wire [7:0] v53; assign v53[7:0] = inp[431:424]; // 0.0
    wire [7:0] v54; assign v54[7:0] = inp[439:432]; // 0.0
    wire [7:0] v55; assign v55[7:0] = inp[447:440]; // 0.0
    wire [7:0] v56; assign v56[7:0] = inp[455:448]; // 0.0
    wire [7:0] v57; assign v57[7:0] = inp[463:456]; // 0.0
    wire [7:0] v58; assign v58[7:0] = inp[471:464]; // 0.0
    wire [7:0] v59; assign v59[7:0] = inp[479:472]; // 0.0
    wire [7:0] v60; assign v60[7:0] = inp[487:480]; // 0.0
    wire [7:0] v61; assign v61[7:0] = inp[495:488]; // 0.0
    wire [7:0] v62; assign v62[7:0] = inp[503:496]; // 0.0
    wire [7:0] v63; assign v63[7:0] = inp[511:504]; // 0.0
    wire [7:0] v64; assign v64[7:0] = v61[7:0]; // 0.0
    wire [7:0] v65; assign v65[7:0] = v2[7:0]; // 0.0
    wire [7:0] v66; assign v66[7:0] = v6[7:0]; // 0.0
    wire [7:0] v67; assign v67[7:0] = v52[7:0]; // 0.0
    wire [7:0] v68; assign v68[7:0] = v56[7:0]; // 0.0
    wire [7:0] v69; assign v69[7:0] = v4[7:0]; // 0.0
    wire [7:0] v70; assign v70[7:0] = v19[7:0]; // 0.0
    wire [7:0] v71; assign v71[7:0] = v62[7:0]; // 0.0
    wire [7:0] v72; assign v72[7:0] = v54[7:0]; // 0.0
    wire [7:0] v73; assign v73[7:0] = v36[7:0]; // 0.0
    wire [7:0] v74; assign v74[7:0] = v32[7:0]; // 0.0
    wire [7:0] v75; assign v75[7:0] = v0[7:0]; // 0.0
    wire [7:0] v76; assign v76[7:0] = v63[7:0]; // 0.0
    wire [7:0] v77; assign v77[7:0] = v59[7:0]; // 0.0
    wire [7:0] v78; assign v78[7:0] = v34[7:0]; // 0.0
    wire [7:0] v79; assign v79[7:0] = v40[7:0]; // 0.0
    wire [7:0] v80; assign v80[7:0] = v41[7:0]; // 0.0
    wire [7:0] v81; assign v81[7:0] = v58[7:0]; // 0.0
    wire [7:0] v82; assign v82[7:0] = v10[7:0]; // 0.0
    wire [7:0] v83; assign v83[7:0] = v33[7:0]; // 0.0
    wire [7:0] v84; assign v84[7:0] = v22[7:0]; // 0.0
    wire [7:0] v85; assign v85[7:0] = v43[7:0]; // 0.0
    wire [7:0] v86; assign v86[7:0] = v49[7:0]; // 0.0
    wire [7:0] v87; assign v87[7:0] = v7[7:0]; // 0.0
    wire [7:0] v88; assign v88[7:0] = v27[7:0]; // 0.0
    wire [7:0] v89; assign v89[7:0] = v44[7:0]; // 0.0
    wire [7:0] v90; assign v90[7:0] = v50[7:0]; // 0.0
    wire [7:0] v91; assign v91[7:0] = v28[7:0]; // 0.0
    wire [7:0] v92; assign v92[7:0] = v48[7:0]; // 0.0
    wire [7:0] v93; assign v93[7:0] = v45[7:0]; // 0.0
    wire [7:0] v94; assign v94[7:0] = v47[7:0]; // 0.0
    wire [7:0] v95; assign v95[7:0] = v21[7:0]; // 0.0
    wire [7:0] v96; assign v96[7:0] = v13[7:0]; // 0.0
    wire [7:0] v97; assign v97[7:0] = v17[7:0]; // 0.0
    wire [7:0] v98; assign v98[7:0] = v38[7:0]; // 0.0
    wire [7:0] v99; assign v99[7:0] = v12[7:0]; // 0.0
    wire [7:0] v100; assign v100[7:0] = v24[7:0]; // 0.0
    wire [7:0] v101; assign v101[7:0] = v23[7:0]; // 0.0
    wire [7:0] v102; assign v102[7:0] = v39[7:0]; // 0.0
    wire [7:0] v103; assign v103[7:0] = v1[7:0]; // 0.0
    wire [7:0] v104; assign v104[7:0] = v15[7:0]; // 0.0
    wire [7:0] v105; assign v105[7:0] = v29[7:0]; // 0.0
    wire [7:0] v106; assign v106[7:0] = v9[7:0]; // 0.0
    wire [7:0] v107; assign v107[7:0] = v51[7:0]; // 0.0
    wire [7:0] v108; assign v108[7:0] = v57[7:0]; // 0.0
    wire [7:0] v109; assign v109[7:0] = v14[7:0]; // 0.0
    wire [7:0] v110; assign v110[7:0] = v42[7:0]; // 0.0
    wire [7:0] v111; assign v111[7:0] = v3[7:0]; // 0.0
    wire [7:0] v112; assign v112[7:0] = v31[7:0]; // 0.0
    wire [7:0] v113; assign v113[7:0] = v60[7:0]; // 0.0
    wire [7:0] v114; assign v114[7:0] = v25[7:0]; // 0.0
    wire [7:0] v115; assign v115[7:0] = v35[7:0]; // 0.0
    wire [7:0] v116; assign v116[7:0] = v30[7:0]; // 0.0
    wire [7:0] v117; assign v117[7:0] = v55[7:0]; // 0.0
    wire [7:0] v118; assign v118[7:0] = v16[7:0]; // 0.0
    wire [7:0] v119; assign v119[7:0] = v20[7:0]; // 0.0
    wire [7:0] v120; assign v120[7:0] = v53[7:0]; // 0.0
    wire [7:0] v121; assign v121[7:0] = v8[7:0]; // 0.0
    wire [7:0] v122; assign v122[7:0] = v37[7:0]; // 0.0
    wire [7:0] v123; assign v123[7:0] = v18[7:0]; // 0.0
    wire [7:0] v124; assign v124[7:0] = v11[7:0]; // 0.0
    wire [7:0] v125; assign v125[7:0] = v46[7:0]; // 0.0
    wire [7:0] v126; assign v126[7:0] = v26[7:0]; // 0.0
    wire [7:0] v127; assign v127[7:0] = v5[7:0]; // 0.0
    wire [8:0] v128; shift_adder #(8, 8, 1, 1, 9, 0, 1) op_128 (v65[7:0], v66[7:0], v128[8:0]); // 1.0
    wire [10:0] v129; shift_adder #(8, 8, 1, 1, 11, 2, 0) op_129 (v67[7:0], v68[7:0], v129[10:0]); // 1.0
    wire [9:0] v130; shift_adder #(8, 8, 1, 1, 10, 1, 0) op_130 (v69[7:0], v70[7:0], v130[9:0]); // 1.0
    wire [10:0] v131; shift_adder #(8, 8, 1, 1, 11, -2, 1) op_131 (v71[7:0], v71[7:0], v131[10:0]); // 1.0
    wire [10:0] v132; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_132 (v73[7:0], v73[7:0], v132[10:0]); // 1.0
    wire [10:0] v133; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_133 (v74[7:0], v74[7:0], v133[10:0]); // 1.0
    wire [10:0] v134; shift_adder #(8, 8, 1, 1, 11, -2, 1) op_134 (v75[7:0], v75[7:0], v134[10:0]); // 1.0
    wire [10:0] v135; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_135 (v76[7:0], v76[7:0], v135[10:0]); // 1.0
    wire [10:0] v136; shift_adder #(8, 8, 1, 1, 11, -2, 1) op_136 (v77[7:0], v77[7:0], v136[10:0]); // 1.0
    wire [11:0] v137; shift_adder #(8, 8, 1, 1, 12, -3, 1) op_137 (v78[7:0], v78[7:0], v137[11:0]); // 1.0
    wire [8:0] v138; shift_adder #(8, 8, 1, 1, 9, 0, 0) op_138 (v79[7:0], v80[7:0], v138[8:0]); // 1.0
    wire [10:0] v139; shift_adder #(8, 8, 1, 1, 11, -2, 1) op_139 (v81[7:0], v81[7:0], v139[10:0]); // 1.0
    wire [10:0] v140; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_140 (v82[7:0], v82[7:0], v140[10:0]); // 1.0
    wire [10:0] v141; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_141 (v83[7:0], v83[7:0], v141[10:0]); // 1.0
    wire [10:0] v142; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_142 (v84[7:0], v84[7:0], v142[10:0]); // 1.0
    wire [16:0] v143; shift_adder #(8, 8, 1, 1, 17, 8, 1) op_143 (v85[7:0], v86[7:0], v143[16:0]); // 1.0
    wire [10:0] v144; shift_adder #(8, 8, 1, 1, 11, -2, 1) op_144 (v80[7:0], v80[7:0], v144[10:0]); // 1.0
    wire [10:0] v145; shift_adder #(8, 8, 1, 1, 11, -2, 1) op_145 (v87[7:0], v87[7:0], v145[10:0]); // 1.0
    wire [11:0] v146; shift_adder #(8, 8, 1, 1, 12, -3, 1) op_146 (v88[7:0], v88[7:0], v146[11:0]); // 1.0
    wire [10:0] v147; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_147 (v89[7:0], v89[7:0], v147[10:0]); // 1.0
    wire [10:0] v148; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_148 (v90[7:0], v90[7:0], v148[10:0]); // 1.0
    wire [12:0] v149; shift_adder #(8, 8, 1, 1, 13, 4, 0) op_149 (v91[7:0], v92[7:0], v149[12:0]); // 1.0
    wire [10:0] v150; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_150 (v93[7:0], v93[7:0], v150[10:0]); // 1.0
    wire [11:0] v151; shift_adder #(8, 8, 1, 1, 12, -3, 0) op_151 (v94[7:0], v94[7:0], v151[11:0]); // 1.0
    wire [10:0] v152; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_152 (v95[7:0], v95[7:0], v152[10:0]); // 1.0
    wire [10:0] v153; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_153 (v96[7:0], v96[7:0], v153[10:0]); // 1.0
    wire [10:0] v154; shift_adder #(8, 8, 1, 1, 11, -2, 1) op_154 (v96[7:0], v96[7:0], v154[10:0]); // 1.0
    wire [10:0] v155; shift_adder #(8, 8, 1, 1, 11, -2, 1) op_155 (v76[7:0], v76[7:0], v155[10:0]); // 1.0
    wire [10:0] v156; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_156 (v97[7:0], v97[7:0], v156[10:0]); // 1.0
    wire [10:0] v157; shift_adder #(8, 8, 1, 1, 11, -2, 1) op_157 (v98[7:0], v98[7:0], v157[10:0]); // 1.0
    wire [10:0] v158; shift_adder #(8, 8, 1, 1, 11, -2, 1) op_158 (v66[7:0], v66[7:0], v158[10:0]); // 1.0
    wire [11:0] v159; shift_adder #(8, 8, 1, 1, 12, -3, 1) op_159 (v99[7:0], v99[7:0], v159[11:0]); // 1.0
    wire [24:0] v160; shift_adder #(8, 8, 1, 1, 25, 16, 0) op_160 (v100[7:0], v101[7:0], v160[24:0]); // 1.0
    wire [10:0] v161; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_161 (v102[7:0], v102[7:0], v161[10:0]); // 1.0
    wire [10:0] v162; shift_adder #(8, 8, 1, 1, 11, -2, 1) op_162 (v69[7:0], v69[7:0], v162[10:0]); // 1.0
    wire [10:0] v163; shift_adder #(8, 8, 1, 1, 11, -2, 1) op_163 (v83[7:0], v83[7:0], v163[10:0]); // 1.0
    wire [11:0] v164; shift_adder #(8, 8, 1, 1, 12, -3, 1) op_164 (v66[7:0], v66[7:0], v164[11:0]); // 1.0
    wire [10:0] v165; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_165 (v103[7:0], v103[7:0], v165[10:0]); // 1.0
    wire [15:0] v166; shift_adder #(8, 8, 1, 1, 16, -7, 0) op_166 (v104[7:0], v80[7:0], v166[15:0]); // 1.0
    wire [17:0] v167; shift_adder #(8, 8, 1, 1, 18, -9, 1) op_167 (v84[7:0], v105[7:0], v167[17:0]); // 1.0
    wire [10:0] v168; shift_adder #(8, 8, 1, 1, 11, -2, 1) op_168 (v65[7:0], v65[7:0], v168[10:0]); // 1.0
    wire [10:0] v169; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_169 (v106[7:0], v106[7:0], v169[10:0]); // 1.0
    wire [9:0] v170; shift_adder #(8, 8, 1, 1, 10, -1, 0) op_170 (v77[7:0], v76[7:0], v170[9:0]); // 1.0
    wire [10:0] v171; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_171 (v107[7:0], v107[7:0], v171[10:0]); // 1.0
    wire [10:0] v172; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_172 (v108[7:0], v108[7:0], v172[10:0]); // 1.0
    wire [10:0] v173; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_173 (v109[7:0], v109[7:0], v173[10:0]); // 1.0
    wire [11:0] v174; shift_adder #(8, 8, 1, 1, 12, 3, 0) op_174 (v91[7:0], v92[7:0], v174[11:0]); // 1.0
    wire [10:0] v175; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_175 (v110[7:0], v110[7:0], v175[10:0]); // 1.0
    wire [10:0] v176; shift_adder #(8, 8, 1, 1, 11, -2, 1) op_176 (v82[7:0], v82[7:0], v176[10:0]); // 1.0
    wire [10:0] v177; shift_adder #(8, 8, 1, 1, 11, -2, 1) op_177 (v111[7:0], v111[7:0], v177[10:0]); // 1.0
    wire [10:0] v178; shift_adder #(8, 8, 1, 1, 11, -2, 1) op_178 (v72[7:0], v72[7:0], v178[10:0]); // 1.0
    wire [10:0] v179; shift_adder #(8, 8, 1, 1, 11, 2, 1) op_179 (v91[7:0], v85[7:0], v179[10:0]); // 1.0
    wire [11:0] v180; shift_adder #(8, 8, 1, 1, 12, -3, 0) op_180 (v81[7:0], v81[7:0], v180[11:0]); // 1.0
    wire [10:0] v181; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_181 (v68[7:0], v68[7:0], v181[10:0]); // 1.0
    wire [10:0] v182; shift_adder #(8, 8, 1, 1, 11, -2, 1) op_182 (v100[7:0], v100[7:0], v182[10:0]); // 1.0
    wire [11:0] v183; shift_adder #(8, 8, 1, 1, 12, -3, 0) op_183 (v74[7:0], v74[7:0], v183[11:0]); // 1.0
    wire [11:0] v184; shift_adder #(8, 8, 1, 1, 12, -3, 0) op_184 (v113[7:0], v113[7:0], v184[11:0]); // 1.0
    wire [10:0] v185; shift_adder #(8, 8, 1, 1, 11, -2, 1) op_185 (v68[7:0], v68[7:0], v185[10:0]); // 1.0
    wire [11:0] v186; shift_adder #(8, 8, 1, 1, 12, 3, 0) op_186 (v102[7:0], v70[7:0], v186[11:0]); // 1.0
    wire [10:0] v187; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_187 (v115[7:0], v115[7:0], v187[10:0]); // 1.0
    wire [10:0] v188; shift_adder #(8, 8, 1, 1, 11, -2, 1) op_188 (v88[7:0], v88[7:0], v188[10:0]); // 1.0
    wire [12:0] v189; shift_adder #(8, 8, 1, 1, 13, -4, 0) op_189 (v114[7:0], v116[7:0], v189[12:0]); // 1.0
    wire [10:0] v190; shift_adder #(8, 8, 1, 1, 11, -2, 1) op_190 (v117[7:0], v117[7:0], v190[10:0]); // 1.0
    wire [10:0] v191; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_191 (v77[7:0], v77[7:0], v191[10:0]); // 1.0
    wire [12:0] v192; shift_adder #(8, 8, 1, 1, 13, -4, 1) op_192 (v105[7:0], v81[7:0], v192[12:0]); // 1.0
    wire [10:0] v193; shift_adder #(8, 8, 1, 1, 11, -2, 1) op_193 (v118[7:0], v118[7:0], v193[10:0]); // 1.0
    wire [11:0] v194; shift_adder #(8, 8, 1, 1, 12, -3, 0) op_194 (v82[7:0], v82[7:0], v194[11:0]); // 1.0
    wire [10:0] v195; shift_adder #(8, 8, 1, 1, 11, -2, 1) op_195 (v85[7:0], v85[7:0], v195[10:0]); // 1.0
    wire [18:0] v196; shift_adder #(8, 8, 1, 1, 19, -10, 0) op_196 (v105[7:0], v110[7:0], v196[18:0]); // 1.0
    wire [10:0] v197; shift_adder #(8, 8, 1, 1, 11, -2, 1) op_197 (v89[7:0], v89[7:0], v197[10:0]); // 1.0
    wire [12:0] v198; shift_adder #(8, 8, 1, 1, 13, 4, 0) op_198 (v66[7:0], v102[7:0], v198[12:0]); // 1.0
    wire [10:0] v199; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_199 (v64[7:0], v64[7:0], v199[10:0]); // 1.0
    wire [10:0] v200; shift_adder #(8, 8, 1, 1, 11, -2, 1) op_200 (v84[7:0], v84[7:0], v200[10:0]); // 1.0
    wire [10:0] v201; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_201 (v119[7:0], v119[7:0], v201[10:0]); // 1.0
    wire [11:0] v202; shift_adder #(8, 8, 1, 1, 12, -3, 0) op_202 (v86[7:0], v86[7:0], v202[11:0]); // 1.0
    wire [10:0] v203; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_203 (v120[7:0], v120[7:0], v203[10:0]); // 1.0
    wire [11:0] v204; shift_adder #(8, 8, 1, 1, 12, -3, 1) op_204 (v73[7:0], v73[7:0], v204[11:0]); // 1.0
    wire [11:0] v205; shift_adder #(8, 8, 1, 1, 12, -3, 1) op_205 (v121[7:0], v121[7:0], v205[11:0]); // 1.0
    wire [10:0] v206; shift_adder #(8, 8, 1, 1, 11, -2, 1) op_206 (v99[7:0], v99[7:0], v206[10:0]); // 1.0
    wire [11:0] v207; shift_adder #(8, 8, 1, 1, 12, -3, 1) op_207 (v69[7:0], v119[7:0], v207[11:0]); // 1.0
    wire [10:0] v208; shift_adder #(8, 8, 1, 1, 11, -2, 1) op_208 (v94[7:0], v94[7:0], v208[10:0]); // 1.0
    wire [10:0] v209; shift_adder #(8, 8, 1, 1, 11, -2, 1) op_209 (v104[7:0], v104[7:0], v209[10:0]); // 1.0
    wire [10:0] v210; shift_adder #(8, 8, 1, 1, 11, -2, 1) op_210 (v105[7:0], v105[7:0], v210[10:0]); // 1.0
    wire [10:0] v211; shift_adder #(8, 8, 1, 1, 11, -2, 1) op_211 (v122[7:0], v122[7:0], v211[10:0]); // 1.0
    wire [10:0] v212; shift_adder #(8, 8, 1, 1, 11, -2, 1) op_212 (v110[7:0], v110[7:0], v212[10:0]); // 1.0
    wire [10:0] v213; shift_adder #(8, 8, 1, 1, 11, -2, 1) op_213 (v67[7:0], v67[7:0], v213[10:0]); // 1.0
    wire [11:0] v214; shift_adder #(8, 8, 1, 1, 12, -3, 0) op_214 (v123[7:0], v123[7:0], v214[11:0]); // 1.0
    wire [10:0] v215; shift_adder #(8, 8, 1, 1, 11, -2, 1) op_215 (v121[7:0], v121[7:0], v215[10:0]); // 1.0
    wire [10:0] v216; shift_adder #(8, 8, 1, 1, 11, -2, 1) op_216 (v116[7:0], v116[7:0], v216[10:0]); // 1.0
    wire [10:0] v217; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_217 (v101[7:0], v101[7:0], v217[10:0]); // 1.0
    wire [10:0] v218; shift_adder #(8, 8, 1, 1, 11, -2, 1) op_218 (v124[7:0], v124[7:0], v218[10:0]); // 1.0
    wire [10:0] v219; shift_adder #(8, 8, 1, 1, 11, -2, 1) op_219 (v123[7:0], v123[7:0], v219[10:0]); // 1.0
    wire [8:0] v220; shift_adder #(8, 8, 1, 1, 9, 0, 1) op_220 (v100[7:0], v92[7:0], v220[8:0]); // 1.0
    wire [8:0] v221; shift_adder #(8, 8, 1, 1, 9, 0, 1) op_221 (v103[7:0], v74[7:0], v221[8:0]); // 1.0
    wire [9:0] v222; shift_adder #(8, 8, 1, 1, 10, 1, 1) op_222 (v87[7:0], v125[7:0], v222[9:0]); // 1.0
    wire [10:0] v223; shift_adder #(8, 8, 1, 1, 11, -2, 1) op_223 (v106[7:0], v106[7:0], v223[10:0]); // 1.0
    wire [11:0] v224; shift_adder #(8, 8, 1, 1, 12, -3, 1) op_224 (v67[7:0], v67[7:0], v224[11:0]); // 1.0
    wire [9:0] v225; shift_adder #(8, 8, 1, 1, 10, 1, 0) op_225 (v97[7:0], v112[7:0], v225[9:0]); // 1.0
    wire [13:0] v226; shift_adder #(8, 8, 1, 1, 14, -5, 1) op_226 (v99[7:0], v117[7:0], v226[13:0]); // 1.0
    wire [11:0] v227; shift_adder #(8, 8, 1, 1, 12, -3, 0) op_227 (v103[7:0], v103[7:0], v227[11:0]); // 1.0
    wire [10:0] v228; shift_adder #(8, 8, 1, 1, 11, -2, 1) op_228 (v114[7:0], v114[7:0], v228[10:0]); // 1.0
    wire [10:0] v229; shift_adder #(8, 8, 1, 1, 11, -2, 1) op_229 (v74[7:0], v74[7:0], v229[10:0]); // 1.0
    wire [8:0] v230; shift_adder #(8, 8, 1, 1, 9, 0, 0) op_230 (v94[7:0], v107[7:0], v230[8:0]); // 1.0
    wire [8:0] v231; shift_adder #(8, 8, 1, 1, 9, 0, 0) op_231 (v123[7:0], v126[7:0], v231[8:0]); // 1.0
    wire [10:0] v232; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_232 (v72[7:0], v72[7:0], v232[10:0]); // 1.0
    wire [10:0] v233; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_233 (v126[7:0], v126[7:0], v233[10:0]); // 1.0
    wire [10:0] v234; shift_adder #(8, 8, 1, 1, 11, -2, 1) op_234 (v101[7:0], v101[7:0], v234[10:0]); // 1.0
    wire [9:0] v235; shift_adder #(8, 8, 1, 1, 10, -1, 0) op_235 (v126[7:0], v91[7:0], v235[9:0]); // 1.0
    wire [13:0] v236; shift_adder #(8, 8, 1, 1, 14, -5, 0) op_236 (v109[7:0], v100[7:0], v236[13:0]); // 1.0
    wire [10:0] v237; shift_adder #(8, 8, 1, 1, 11, -2, 1) op_237 (v79[7:0], v79[7:0], v237[10:0]); // 1.0
    wire [10:0] v238; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_238 (v65[7:0], v65[7:0], v238[10:0]); // 1.0
    wire [11:0] v239; shift_adder #(8, 8, 1, 1, 12, 3, 0) op_239 (v126[7:0], v91[7:0], v239[11:0]); // 1.0
    wire [15:0] v240; shift_adder #(8, 8, 1, 1, 16, 7, 1) op_240 (v65[7:0], v97[7:0], v240[15:0]); // 1.0
    wire [10:0] v241; shift_adder #(8, 8, 1, 1, 11, -2, 1) op_241 (v127[7:0], v127[7:0], v241[10:0]); // 1.0
    wire [10:0] v242; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_242 (v111[7:0], v111[7:0], v242[10:0]); // 1.0
    wire [11:0] v243; shift_adder #(8, 8, 1, 1, 12, -3, 0) op_243 (v122[7:0], v122[7:0], v243[11:0]); // 1.0
    wire [10:0] v244; shift_adder #(8, 8, 1, 1, 11, -2, 1) op_244 (v112[7:0], v112[7:0], v244[10:0]); // 1.0
    wire [10:0] v245; shift_adder #(8, 8, 1, 1, 11, -2, 1) op_245 (v126[7:0], v126[7:0], v245[10:0]); // 1.0
    wire [10:0] v246; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_246 (v113[7:0], v113[7:0], v246[10:0]); // 1.0
    wire [11:0] v247; shift_adder #(8, 8, 1, 1, 12, -3, 0) op_247 (v75[7:0], v75[7:0], v247[11:0]); // 1.0
    wire [9:0] v248; shift_adder #(8, 8, 1, 1, 10, 1, 0) op_248 (v104[7:0], v116[7:0], v248[9:0]); // 1.0
    wire [13:0] v249; shift_adder #(8, 8, 1, 1, 14, -5, 1) op_249 (v121[7:0], v68[7:0], v249[13:0]); // 1.0
    wire [10:0] v250; shift_adder #(8, 8, 1, 1, 11, -2, 1) op_250 (v119[7:0], v119[7:0], v250[10:0]); // 1.0
    wire [10:0] v251; shift_adder #(8, 8, 1, 1, 11, -2, 1) op_251 (v93[7:0], v93[7:0], v251[10:0]); // 1.0
    wire [9:0] v252; shift_adder #(8, 8, 1, 1, 10, 1, 0) op_252 (v82[7:0], v91[7:0], v252[9:0]); // 1.0
    wire [14:0] v253; shift_adder #(8, 8, 1, 1, 15, -6, 0) op_253 (v127[7:0], v120[7:0], v253[14:0]); // 1.0
    wire [9:0] v254; shift_adder #(8, 8, 1, 1, 10, -1, 0) op_254 (v115[7:0], v117[7:0], v254[9:0]); // 1.0
    wire [10:0] v255; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_255 (v98[7:0], v98[7:0], v255[10:0]); // 1.0
    wire [8:0] v256; shift_adder #(8, 8, 1, 1, 9, 0, 1) op_256 (v104[7:0], v80[7:0], v256[8:0]); // 1.0
    wire [11:0] v257; shift_adder #(8, 8, 1, 1, 12, -3, 0) op_257 (v96[7:0], v96[7:0], v257[11:0]); // 1.0
    wire [22:0] v258; shift_adder #(8, 8, 1, 1, 23, -14, 1) op_258 (v115[7:0], v102[7:0], v258[22:0]); // 1.0
    wire [10:0] v259; shift_adder #(8, 8, 1, 1, 11, -2, 1) op_259 (v78[7:0], v78[7:0], v259[10:0]); // 1.0
    wire [9:0] v260; shift_adder #(8, 8, 1, 1, 10, 1, 1) op_260 (v109[7:0], v117[7:0], v260[9:0]); // 1.0
    wire [24:0] v261; shift_adder #(8, 8, 1, 1, 25, -16, 1) op_261 (v88[7:0], v88[7:0], v261[24:0]); // 1.0
    wire [31:0] v262; shift_adder #(8, 8, 1, 1, 32, -23, 1) op_262 (v89[7:0], v96[7:0], v262[31:0]); // 1.0
    wire [9:0] v263; shift_adder #(8, 8, 1, 1, 10, -1, 1) op_263 (v119[7:0], v101[7:0], v263[9:0]); // 1.0
    wire [10:0] v264; shift_adder #(8, 8, 1, 1, 11, -2, 1) op_264 (v70[7:0], v70[7:0], v264[10:0]); // 1.0
    wire [11:0] v265; shift_adder #(8, 8, 1, 1, 12, -3, 0) op_265 (v98[7:0], v98[7:0], v265[11:0]); // 1.0
    wire [10:0] v266; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_266 (v79[7:0], v79[7:0], v266[10:0]); // 1.0
    wire [11:0] v267; shift_adder #(8, 8, 1, 1, 12, -3, 1) op_267 (v88[7:0], v92[7:0], v267[11:0]); // 1.0
    wire [10:0] v268; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_268 (v116[7:0], v116[7:0], v268[10:0]); // 1.0
    wire [10:0] v269; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_269 (v100[7:0], v100[7:0], v269[10:0]); // 1.0
    wire [10:0] v270; shift_adder #(8, 8, 1, 1, 11, -2, 1) op_270 (v86[7:0], v86[7:0], v270[10:0]); // 1.0
    wire [13:0] v271; shift_adder #(8, 8, 1, 1, 14, -5, 1) op_271 (v97[7:0], v64[7:0], v271[13:0]); // 1.0
    wire [12:0] v272; shift_adder #(8, 8, 1, 1, 13, 4, 0) op_272 (v83[7:0], v73[7:0], v272[12:0]); // 1.0
    wire [9:0] v273; shift_adder #(8, 8, 1, 1, 10, 1, 0) op_273 (v70[7:0], v83[7:0], v273[9:0]); // 1.0
    wire [10:0] v274; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_274 (v95[7:0], v85[7:0], v274[10:0]); // 1.0
    wire [10:0] v275; shift_adder #(8, 8, 1, 1, 11, -2, 1) op_275 (v113[7:0], v113[7:0], v275[10:0]); // 1.0
    wire [10:0] v276; shift_adder #(8, 8, 1, 1, 11, -2, 1) op_276 (v125[7:0], v125[7:0], v276[10:0]); // 1.0
    wire [10:0] v277; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_277 (v123[7:0], v123[7:0], v277[10:0]); // 1.0
    wire [12:0] v278; shift_adder #(8, 8, 1, 1, 13, -4, 0) op_278 (v102[7:0], v103[7:0], v278[12:0]); // 1.0
    wire [11:0] v279; shift_adder #(8, 8, 1, 1, 12, -3, 1) op_279 (v125[7:0], v90[7:0], v279[11:0]); // 1.0
    wire [11:0] v280; shift_adder #(8, 8, 1, 1, 12, -3, 1) op_280 (v109[7:0], v109[7:0], v280[11:0]); // 1.0
    wire [10:0] v281; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_281 (v87[7:0], v124[7:0], v281[10:0]); // 1.0
    wire [9:0] v282; shift_adder #(8, 8, 1, 1, 10, 1, 1) op_282 (v104[7:0], v79[7:0], v282[9:0]); // 1.0
    wire [10:0] v283; shift_adder #(8, 8, 1, 1, 11, -2, 1) op_283 (v115[7:0], v115[7:0], v283[10:0]); // 1.0
    wire [10:0] v284; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_284 (v117[7:0], v117[7:0], v284[10:0]); // 1.0
    wire [11:0] v285; shift_adder #(8, 8, 1, 1, 12, 3, 0) op_285 (v87[7:0], v125[7:0], v285[11:0]); // 1.0
    wire [17:0] v286; shift_adder #(8, 8, 1, 1, 18, -9, 1) op_286 (v97[7:0], v71[7:0], v286[17:0]); // 1.0
    wire [10:0] v287; shift_adder #(8, 8, 1, 1, 11, 2, 1) op_287 (v91[7:0], v92[7:0], v287[10:0]); // 1.0
    wire [11:0] v288; shift_adder #(8, 8, 1, 1, 12, -3, 0) op_288 (v70[7:0], v70[7:0], v288[11:0]); // 1.0
    wire [10:0] v289; shift_adder #(8, 8, 1, 1, 11, -2, 1) op_289 (v95[7:0], v95[7:0], v289[10:0]); // 1.0
    wire [13:0] v290; shift_adder #(8, 8, 1, 1, 14, 5, 0) op_290 (v127[7:0], v106[7:0], v290[13:0]); // 1.0
    wire [9:0] v291; shift_adder #(8, 8, 1, 1, 10, -1, 0) op_291 (v96[7:0], v89[7:0], v291[9:0]); // 1.0
    wire [11:0] v292; shift_adder #(8, 8, 1, 1, 12, 3, 1) op_292 (v91[7:0], v92[7:0], v292[11:0]); // 1.0
    wire [10:0] v293; shift_adder #(8, 8, 1, 1, 11, -2, 1) op_293 (v90[7:0], v90[7:0], v293[10:0]); // 1.0
    wire [10:0] v294; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_294 (v78[7:0], v78[7:0], v294[10:0]); // 1.0
    wire [14:0] v295; shift_adder #(8, 8, 1, 1, 15, 6, 1) op_295 (v127[7:0], v108[7:0], v295[14:0]); // 1.0
    wire [12:0] v296; shift_adder #(8, 8, 1, 1, 13, -4, 0) op_296 (v114[7:0], v114[7:0], v296[12:0]); // 1.0
    wire [10:0] v297; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_297 (v75[7:0], v75[7:0], v297[10:0]); // 1.0
    wire [10:0] v298; shift_adder #(8, 8, 1, 1, 11, -2, 1) op_298 (v97[7:0], v97[7:0], v298[10:0]); // 1.0
    wire [10:0] v299; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_299 (v114[7:0], v114[7:0], v299[10:0]); // 1.0
    wire [10:0] v300; shift_adder #(8, 8, 1, 1, 11, -2, 1) op_300 (v120[7:0], v120[7:0], v300[10:0]); // 1.0
    wire [10:0] v301; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_301 (v88[7:0], v88[7:0], v301[10:0]); // 1.0
    wire [8:0] v302; shift_adder #(8, 8, 1, 1, 9, 0, 0) op_302 (v111[7:0], v66[7:0], v302[8:0]); // 1.0
    wire [10:0] v303; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_303 (v94[7:0], v94[7:0], v303[10:0]); // 1.0
    wire [11:0] v304; shift_adder #(8, 8, 1, 1, 12, -3, 0) op_304 (v65[7:0], v65[7:0], v304[11:0]); // 1.0
    wire [11:0] v305; shift_adder #(8, 8, 1, 1, 12, -3, 0) op_305 (v108[7:0], v108[7:0], v305[11:0]); // 1.0
    wire [16:0] v306; shift_adder #(8, 8, 1, 1, 17, -8, 0) op_306 (v74[7:0], v108[7:0], v306[16:0]); // 1.0
    wire [9:0] v307; shift_adder #(8, 8, 1, 1, 10, 1, 1) op_307 (v122[7:0], v113[7:0], v307[9:0]); // 1.0
    wire [14:0] v308; shift_adder #(8, 8, 1, 1, 15, 6, 1) op_308 (v106[7:0], v125[7:0], v308[14:0]); // 1.0
    wire [8:0] v309; shift_adder #(8, 8, 1, 1, 9, 0, 0) op_309 (v121[7:0], v114[7:0], v309[8:0]); // 1.0
    wire [19:0] v310; shift_adder #(8, 8, 1, 1, 20, -11, 1) op_310 (v81[7:0], v76[7:0], v310[19:0]); // 1.0
    wire [9:0] v311; shift_adder #(8, 8, 1, 1, 10, 1, 1) op_311 (v101[7:0], v100[7:0], v311[9:0]); // 1.0
    wire [10:0] v312; shift_adder #(8, 8, 1, 1, 11, 2, 0) op_312 (v106[7:0], v73[7:0], v312[10:0]); // 1.0
    wire [14:0] v313; shift_adder #(8, 8, 1, 1, 15, -6, 1) op_313 (v104[7:0], v108[7:0], v313[14:0]); // 1.0
    wire [11:0] v314; shift_adder #(8, 8, 1, 1, 12, -3, 0) op_314 (v111[7:0], v111[7:0], v314[11:0]); // 1.0
    wire [18:0] v315; shift_adder #(8, 8, 1, 1, 19, 10, 0) op_315 (v82[7:0], v93[7:0], v315[18:0]); // 1.0
    wire [8:0] v316; shift_adder #(8, 8, 1, 1, 9, 0, 1) op_316 (v95[7:0], v126[7:0], v316[8:0]); // 1.0
    wire [10:0] v317; shift_adder #(8, 8, 1, 1, 11, -2, 1) op_317 (v103[7:0], v103[7:0], v317[10:0]); // 1.0
    wire [14:0] v318; shift_adder #(8, 8, 1, 1, 15, -6, 0) op_318 (v83[7:0], v80[7:0], v318[14:0]); // 1.0
    wire [10:0] v319; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_319 (v104[7:0], v104[7:0], v319[10:0]); // 1.0
    wire [10:0] v320; shift_adder #(8, 8, 1, 1, 11, -2, 1) op_320 (v108[7:0], v108[7:0], v320[10:0]); // 1.0
    wire [11:0] v321; shift_adder #(8, 8, 1, 1, 12, -3, 1) op_321 (v118[7:0], v118[7:0], v321[11:0]); // 1.0
    wire [8:0] v322; shift_adder #(8, 8, 1, 1, 9, 0, 1) op_322 (v107[7:0], v64[7:0], v322[8:0]); // 1.0
    wire [10:0] v323; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_323 (v80[7:0], v80[7:0], v323[10:0]); // 1.0
    wire [10:0] v324; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_324 (v99[7:0], v99[7:0], v324[10:0]); // 1.0
    wire [11:0] v325; shift_adder #(8, 8, 1, 1, 12, 3, 1) op_325 (v84[7:0], v79[7:0], v325[11:0]); // 1.0
    wire [12:0] v326; shift_adder #(8, 8, 1, 1, 13, 4, 0) op_326 (v69[7:0], v110[7:0], v326[12:0]); // 1.0
    wire [12:0] v327; shift_adder #(8, 8, 1, 1, 13, -4, 0) op_327 (v103[7:0], v96[7:0], v327[12:0]); // 1.0
    wire [10:0] v328; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_328 (v127[7:0], v127[7:0], v328[10:0]); // 1.0
    wire [10:0] v329; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_329 (v87[7:0], v87[7:0], v329[10:0]); // 1.0
    wire [10:0] v330; shift_adder #(8, 8, 1, 1, 11, 2, 1) op_330 (v124[7:0], v71[7:0], v330[10:0]); // 1.0
    wire [9:0] v331; shift_adder #(8, 8, 1, 1, 10, 1, 0) op_331 (v115[7:0], v77[7:0], v331[9:0]); // 1.0
    wire [31:0] v332; shift_adder #(8, 8, 1, 1, 32, -23, 1) op_332 (v64[7:0], v83[7:0], v332[31:0]); // 1.0
    wire [11:0] v333; shift_adder #(8, 8, 1, 1, 12, -3, 1) op_333 (v96[7:0], v96[7:0], v333[11:0]); // 1.0
    wire [10:0] v334; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_334 (v66[7:0], v66[7:0], v334[10:0]); // 1.0
    wire [16:0] v335; shift_adder #(8, 8, 1, 1, 17, -8, 1) op_335 (v118[7:0], v85[7:0], v335[16:0]); // 1.0
    wire [11:0] v336; shift_adder #(8, 8, 1, 1, 12, -3, 0) op_336 (v112[7:0], v112[7:0], v336[11:0]); // 1.0
    wire [11:0] v337; shift_adder #(8, 8, 1, 1, 12, -3, 0) op_337 (v76[7:0], v76[7:0], v337[11:0]); // 1.0
    wire [10:0] v338; shift_adder #(8, 8, 1, 1, 11, -2, 1) op_338 (v102[7:0], v102[7:0], v338[10:0]); // 1.0
    wire [11:0] v339; shift_adder #(8, 8, 1, 1, 12, 3, 1) op_339 (v123[7:0], v68[7:0], v339[11:0]); // 1.0
    wire [8:0] v340; shift_adder #(8, 8, 1, 1, 9, 0, 0) op_340 (v75[7:0], v72[7:0], v340[8:0]); // 1.0
    wire [10:0] v341; shift_adder #(8, 8, 1, 1, 11, -2, 1) op_341 (v109[7:0], v109[7:0], v341[10:0]); // 1.0
    wire [13:0] v342; shift_adder #(8, 8, 1, 1, 14, -5, 1) op_342 (v95[7:0], v112[7:0], v342[13:0]); // 1.0
    wire [10:0] v343; shift_adder #(8, 8, 1, 1, 11, 2, 1) op_343 (v69[7:0], v90[7:0], v343[10:0]); // 1.0
    wire [12:0] v344; shift_adder #(8, 8, 1, 1, 13, -4, 0) op_344 (v127[7:0], v124[7:0], v344[12:0]); // 1.0
    wire [10:0] v345; shift_adder #(8, 8, 1, 1, 11, -2, 1) op_345 (v126[7:0], v71[7:0], v345[10:0]); // 1.0
    wire [12:0] v346; shift_adder #(8, 8, 1, 1, 13, -4, 0) op_346 (v78[7:0], v117[7:0], v346[12:0]); // 1.0
    wire [11:0] v347; shift_adder #(8, 8, 1, 1, 12, -3, 1) op_347 (v110[7:0], v110[7:0], v347[11:0]); // 1.0
    wire [16:0] v348; shift_adder #(8, 8, 1, 1, 17, 8, 1) op_348 (v127[7:0], v112[7:0], v348[16:0]); // 1.0
    wire [12:0] v349; shift_adder #(8, 8, 1, 1, 13, -4, 0) op_349 (v117[7:0], v96[7:0], v349[12:0]); // 1.0
    wire [15:0] v350; shift_adder #(8, 8, 1, 1, 16, 7, 1) op_350 (v112[7:0], v94[7:0], v350[15:0]); // 1.0
    wire [8:0] v351; shift_adder #(8, 8, 1, 1, 9, 0, 1) op_351 (v116[7:0], v80[7:0], v351[8:0]); // 1.0
    wire [10:0] v352; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_352 (v81[7:0], v81[7:0], v352[10:0]); // 1.0
    wire [10:0] v353; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_353 (v112[7:0], v112[7:0], v353[10:0]); // 1.0
    wire [11:0] v354; shift_adder #(8, 8, 1, 1, 12, -3, 0) op_354 (v105[7:0], v72[7:0], v354[11:0]); // 1.0
    wire [11:0] v355; shift_adder #(8, 8, 1, 1, 12, 3, 0) op_355 (v114[7:0], v78[7:0], v355[11:0]); // 1.0
    wire [13:0] v356; shift_adder #(8, 8, 1, 1, 14, -5, 0) op_356 (v127[7:0], v74[7:0], v356[13:0]); // 1.0
    wire [11:0] v357; shift_adder #(8, 8, 1, 1, 12, -3, 0) op_357 (v67[7:0], v67[7:0], v357[11:0]); // 1.0
    wire [10:0] v358; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_358 (v105[7:0], v105[7:0], v358[10:0]); // 1.0
    wire [12:0] v359; shift_adder #(8, 8, 1, 1, 13, 4, 1) op_359 (v109[7:0], v79[7:0], v359[12:0]); // 1.0
    wire [8:0] v360; shift_adder #(8, 8, 1, 1, 9, 0, 1) op_360 (v91[7:0], v72[7:0], v360[8:0]); // 1.0
    wire [10:0] v361; shift_adder #(8, 8, 1, 1, 11, -2, 1) op_361 (v73[7:0], v73[7:0], v361[10:0]); // 1.0
    wire [10:0] v362; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_362 (v67[7:0], v67[7:0], v362[10:0]); // 1.0
    wire [11:0] v363; shift_adder #(8, 8, 1, 1, 12, -3, 1) op_363 (v107[7:0], v107[7:0], v363[11:0]); // 1.0
    wire [20:0] v364; shift_adder #(8, 8, 1, 1, 21, -12, 1) op_364 (v109[7:0], v93[7:0], v364[20:0]); // 1.0
    wire [11:0] v365; shift_adder #(8, 8, 1, 1, 12, -3, 1) op_365 (v64[7:0], v64[7:0], v365[11:0]); // 1.0
    wire [9:0] v366; shift_adder #(8, 8, 1, 1, 10, 1, 0) op_366 (v87[7:0], v105[7:0], v366[9:0]); // 1.0
    wire [10:0] v367; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_367 (v125[7:0], v125[7:0], v367[10:0]); // 1.0
    wire [8:0] v368; shift_adder #(8, 8, 1, 1, 9, 0, 0) op_368 (v69[7:0], v115[7:0], v368[8:0]); // 1.0
    wire [8:0] v369; shift_adder #(8, 8, 1, 1, 9, 0, 1) op_369 (v70[7:0], v84[7:0], v369[8:0]); // 1.0
    wire [8:0] v370; shift_adder #(8, 8, 1, 1, 9, 0, 1) op_370 (v96[7:0], v98[7:0], v370[8:0]); // 1.0
    wire [21:0] v371; shift_adder #(8, 8, 1, 1, 22, -13, 1) op_371 (v103[7:0], v127[7:0], v371[21:0]); // 1.0
    wire [11:0] v372; shift_adder #(8, 8, 1, 1, 12, -3, 0) op_372 (v77[7:0], v77[7:0], v372[11:0]); // 1.0
    wire [25:0] v373; shift_adder #(8, 8, 1, 1, 26, -17, 1) op_373 (v119[7:0], v92[7:0], v373[25:0]); // 1.0
    wire [10:0] v374; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_374 (v122[7:0], v122[7:0], v374[10:0]); // 1.0
    wire [10:0] v375; shift_adder #(8, 8, 1, 1, 11, -2, 1) op_375 (v64[7:0], v64[7:0], v375[10:0]); // 1.0
    wire [18:0] v376; shift_adder #(8, 8, 1, 1, 19, 10, 1) op_376 (v85[7:0], v89[7:0], v376[18:0]); // 1.0
    wire [10:0] v377; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_377 (v120[7:0], v113[7:0], v377[10:0]); // 1.0
    wire [17:0] v378; shift_adder #(8, 8, 1, 1, 18, 9, 0) op_378 (v97[7:0], v104[7:0], v378[17:0]); // 1.0
    wire [10:0] v379; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_379 (v70[7:0], v70[7:0], v379[10:0]); // 1.0
    wire [11:0] v380; shift_adder #(8, 8, 1, 1, 12, -3, 0) op_380 (v87[7:0], v87[7:0], v380[11:0]); // 1.0
    wire [30:0] v381; shift_adder #(8, 8, 1, 1, 31, -22, 0) op_381 (v99[7:0], v100[7:0], v381[30:0]); // 1.0
    wire [11:0] v382; shift_adder #(8, 8, 1, 1, 12, -3, 1) op_382 (v68[7:0], v68[7:0], v382[11:0]); // 1.0
    wire [11:0] v383; shift_adder #(8, 8, 1, 1, 12, -3, 0) op_383 (v121[7:0], v121[7:0], v383[11:0]); // 1.0
    wire [8:0] v384; shift_adder #(8, 8, 1, 1, 9, 0, 1) op_384 (v82[7:0], v70[7:0], v384[8:0]); // 1.0
    wire [11:0] v385; shift_adder #(8, 8, 1, 1, 12, -3, 1) op_385 (v108[7:0], v108[7:0], v385[11:0]); // 1.0
    wire [10:0] v386; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_386 (v86[7:0], v86[7:0], v386[10:0]); // 1.0
    wire [11:0] v387; shift_adder #(8, 8, 1, 1, 12, -3, 1) op_387 (v122[7:0], v122[7:0], v387[11:0]); // 1.0
    wire [11:0] v388; shift_adder #(8, 8, 1, 1, 12, -3, 0) op_388 (v105[7:0], v67[7:0], v388[11:0]); // 1.0
    wire [11:0] v389; shift_adder #(8, 8, 1, 1, 12, -3, 0) op_389 (v96[7:0], v89[7:0], v389[11:0]); // 1.0
    wire [15:0] v390; shift_adder #(8, 8, 1, 1, 16, -7, 0) op_390 (v102[7:0], v102[7:0], v390[15:0]); // 1.0
    wire [12:0] v391; shift_adder #(8, 8, 1, 1, 13, 4, 0) op_391 (v98[7:0], v108[7:0], v391[12:0]); // 1.0
    wire [11:0] v392; shift_adder #(8, 8, 1, 1, 12, -3, 1) op_392 (v93[7:0], v93[7:0], v392[11:0]); // 1.0
    wire [10:0] v393; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_393 (v121[7:0], v121[7:0], v393[10:0]); // 1.0
    wire [13:0] v394; shift_adder #(8, 8, 1, 1, 14, -5, 0) op_394 (v119[7:0], v98[7:0], v394[13:0]); // 1.0
    wire [8:0] v395; shift_adder #(8, 8, 1, 1, 9, 0, 0) op_395 (v102[7:0], v117[7:0], v395[8:0]); // 1.0
    wire [10:0] v396; shift_adder #(8, 8, 1, 1, 11, -2, 1) op_396 (v107[7:0], v107[7:0], v396[10:0]); // 1.0
    wire [11:0] v397; shift_adder #(8, 8, 1, 1, 12, -3, 1) op_397 (v85[7:0], v85[7:0], v397[11:0]); // 1.0
    wire [11:0] v398; shift_adder #(8, 8, 1, 1, 12, -3, 1) op_398 (v95[7:0], v95[7:0], v398[11:0]); // 1.0
    wire [33:0] v399; shift_adder #(8, 8, 1, 1, 34, 25, 1) op_399 (v87[7:0], v112[7:0], v399[33:0]); // 1.0
    wire [10:0] v400; shift_adder #(8, 8, 1, 1, 11, 2, 0) op_400 (v103[7:0], v80[7:0], v400[10:0]); // 1.0
    wire [8:0] v401; shift_adder #(8, 8, 1, 1, 9, 0, 0) op_401 (v119[7:0], v72[7:0], v401[8:0]); // 1.0
    wire [11:0] v402; shift_adder #(8, 8, 1, 1, 12, 3, 1) op_402 (v83[7:0], v107[7:0], v402[11:0]); // 1.0
    wire [8:0] v403; shift_adder #(8, 8, 1, 1, 9, 0, 0) op_403 (v97[7:0], v64[7:0], v403[8:0]); // 1.0
    wire [11:0] v404; shift_adder #(8, 8, 1, 1, 12, -3, 1) op_404 (v89[7:0], v94[7:0], v404[11:0]); // 1.0
    wire [8:0] v405; shift_adder #(8, 8, 1, 1, 9, 0, 1) op_405 (v78[7:0], v120[7:0], v405[8:0]); // 1.0
    wire [12:0] v406; shift_adder #(8, 8, 1, 1, 13, -4, 0) op_406 (v87[7:0], v109[7:0], v406[12:0]); // 1.0
    wire [11:0] v407; shift_adder #(8, 8, 1, 1, 12, 3, 1) op_407 (v81[7:0], v76[7:0], v407[11:0]); // 1.0
    wire [11:0] v408; shift_adder #(8, 8, 1, 1, 12, -3, 1) op_408 (v126[7:0], v126[7:0], v408[11:0]); // 1.0
    wire [11:0] v409; shift_adder #(8, 8, 1, 1, 12, -3, 0) op_409 (v99[7:0], v99[7:0], v409[11:0]); // 1.0
    wire [13:0] v410; shift_adder #(8, 8, 1, 1, 14, -5, 1) op_410 (v112[7:0], v125[7:0], v410[13:0]); // 1.0
    wire [11:0] v411; shift_adder #(8, 8, 1, 1, 12, 3, 1) op_411 (v92[7:0], v117[7:0], v411[11:0]); // 1.0
    wire [13:0] v412; shift_adder #(8, 8, 1, 1, 14, 5, 1) op_412 (v114[7:0], v74[7:0], v412[13:0]); // 1.0
    wire [10:0] v413; shift_adder #(8, 8, 1, 1, 11, -2, 1) op_413 (v116[7:0], v93[7:0], v413[10:0]); // 1.0
    wire [16:0] v414; shift_adder #(8, 8, 1, 1, 17, -8, 1) op_414 (v66[7:0], v99[7:0], v414[16:0]); // 1.0
    wire [10:0] v415; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_415 (v82[7:0], v118[7:0], v415[10:0]); // 1.0
    wire [12:0] v416; shift_adder #(8, 8, 1, 1, 13, -4, 1) op_416 (v105[7:0], v71[7:0], v416[12:0]); // 1.0
    wire [13:0] v417; shift_adder #(8, 8, 1, 1, 14, -5, 0) op_417 (v101[7:0], v91[7:0], v417[13:0]); // 1.0
    wire [10:0] v418; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_418 (v69[7:0], v69[7:0], v418[10:0]); // 1.0
    wire [9:0] v419; shift_adder #(8, 8, 1, 1, 10, 1, 0) op_419 (v109[7:0], v116[7:0], v419[9:0]); // 1.0
    wire [10:0] v420; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_420 (v71[7:0], v71[7:0], v420[10:0]); // 1.0
    wire [9:0] v421; shift_adder #(8, 8, 1, 1, 10, 1, 0) op_421 (v86[7:0], v67[7:0], v421[9:0]); // 1.0
    wire [13:0] v422; shift_adder #(8, 8, 1, 1, 14, 5, 0) op_422 (v125[7:0], v83[7:0], v422[13:0]); // 1.0
    wire [11:0] v423; shift_adder #(8, 8, 1, 1, 12, 3, 0) op_423 (v75[7:0], v79[7:0], v423[11:0]); // 1.0
    wire [10:0] v424; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_424 (v96[7:0], v120[7:0], v424[10:0]); // 1.0
    wire [10:0] v425; shift_adder #(8, 8, 1, 1, 11, 2, 0) op_425 (v91[7:0], v92[7:0], v425[10:0]); // 1.0
    wire [15:0] v426; shift_adder #(8, 8, 1, 1, 16, 7, 1) op_426 (v123[7:0], v125[7:0], v426[15:0]); // 1.0
    wire [20:0] v427; shift_adder #(8, 8, 1, 1, 21, -12, 0) op_427 (v93[7:0], v77[7:0], v427[20:0]); // 1.0
    wire [9:0] v428; shift_adder #(8, 8, 1, 1, 10, -1, 0) op_428 (v92[7:0], v76[7:0], v428[9:0]); // 1.0
    wire [17:0] v429; shift_adder #(8, 8, 1, 1, 18, 9, 0) op_429 (v100[7:0], v103[7:0], v429[17:0]); // 1.0
    wire [10:0] v430; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_430 (v124[7:0], v124[7:0], v430[10:0]); // 1.0
    wire [14:0] v431; shift_adder #(8, 8, 1, 1, 15, -6, 1) op_431 (v97[7:0], v93[7:0], v431[14:0]); // 1.0
    wire [9:0] v432; shift_adder #(8, 8, 1, 1, 10, 1, 0) op_432 (v95[7:0], v112[7:0], v432[9:0]); // 1.0
    wire [8:0] v433; shift_adder #(8, 8, 1, 1, 9, 0, 0) op_433 (v127[7:0], v68[7:0], v433[8:0]); // 1.0
    wire [11:0] v434; shift_adder #(8, 8, 1, 1, 12, -3, 1) op_434 (v82[7:0], v82[7:0], v434[11:0]); // 1.0
    wire [9:0] v435; shift_adder #(8, 8, 1, 1, 10, -1, 1) op_435 (v65[7:0], v72[7:0], v435[9:0]); // 1.0
    wire [16:0] v436; shift_adder #(8, 8, 1, 1, 17, 8, 0) op_436 (v104[7:0], v100[7:0], v436[16:0]); // 1.0
    wire [9:0] v437; shift_adder #(8, 8, 1, 1, 10, 1, 0) op_437 (v115[7:0], v98[7:0], v437[9:0]); // 1.0
    wire [11:0] v438; shift_adder #(8, 8, 1, 1, 12, -3, 1) op_438 (v84[7:0], v102[7:0], v438[11:0]); // 1.0
    wire [28:0] v439; shift_adder #(8, 8, 1, 1, 29, -20, 0) op_439 (v70[7:0], v94[7:0], v439[28:0]); // 1.0
    wire [22:0] v440; shift_adder #(8, 8, 1, 1, 23, 14, 0) op_440 (v118[7:0], v100[7:0], v440[22:0]); // 1.0
    wire [8:0] v441; shift_adder #(8, 8, 1, 1, 9, 0, 0) op_441 (v106[7:0], v118[7:0], v441[8:0]); // 1.0
    wire [9:0] v442; shift_adder #(8, 8, 1, 1, 10, 1, 0) op_442 (v104[7:0], v107[7:0], v442[9:0]); // 1.0
    wire [10:0] v443; shift_adder #(8, 8, 1, 1, 11, 2, 0) op_443 (v81[7:0], v71[7:0], v443[10:0]); // 1.0
    wire [13:0] v444; shift_adder #(8, 8, 1, 1, 14, -5, 1) op_444 (v70[7:0], v110[7:0], v444[13:0]); // 1.0
    wire [9:0] v445; shift_adder #(8, 8, 1, 1, 10, 1, 0) op_445 (v97[7:0], v116[7:0], v445[9:0]); // 1.0
    wire [9:0] v446; shift_adder #(8, 8, 1, 1, 10, 1, 0) op_446 (v121[7:0], v125[7:0], v446[9:0]); // 1.0
    wire [11:0] v447; shift_adder #(8, 8, 1, 1, 12, -3, 1) op_447 (v113[7:0], v113[7:0], v447[11:0]); // 1.0
    wire [31:0] v448; shift_adder #(8, 8, 1, 1, 32, -23, 0) op_448 (v74[7:0], v64[7:0], v448[31:0]); // 1.0
    wire [12:0] v449; shift_adder #(8, 8, 1, 1, 13, 4, 0) op_449 (v88[7:0], v64[7:0], v449[12:0]); // 1.0
    wire [9:0] v450; shift_adder #(8, 8, 1, 1, 10, 1, 0) op_450 (v106[7:0], v98[7:0], v450[9:0]); // 1.0
    wire [12:0] v451; shift_adder #(8, 8, 1, 1, 13, 4, 1) op_451 (v95[7:0], v91[7:0], v451[12:0]); // 1.0
    wire [11:0] v452; shift_adder #(8, 8, 1, 1, 12, -3, 0) op_452 (v84[7:0], v84[7:0], v452[11:0]); // 1.0
    wire [11:0] v453; shift_adder #(8, 8, 1, 1, 12, -3, 0) op_453 (v97[7:0], v97[7:0], v453[11:0]); // 1.0
    wire [13:0] v454; shift_adder #(8, 8, 1, 1, 14, -5, 0) op_454 (v94[7:0], v117[7:0], v454[13:0]); // 1.0
    wire [10:0] v455; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_455 (v118[7:0], v118[7:0], v455[10:0]); // 1.0
    wire [14:0] v456; shift_adder #(8, 8, 1, 1, 15, 6, 1) op_456 (v100[7:0], v94[7:0], v456[14:0]); // 1.0
    wire [11:0] v457; shift_adder #(8, 8, 1, 1, 12, -3, 0) op_457 (v83[7:0], v83[7:0], v457[11:0]); // 1.0
    wire [12:0] v458; shift_adder #(8, 8, 1, 1, 13, -4, 1) op_458 (v111[7:0], v81[7:0], v458[12:0]); // 1.0
    wire [9:0] v459; shift_adder #(8, 8, 1, 1, 10, -1, 1) op_459 (v78[7:0], v81[7:0], v459[9:0]); // 1.0
    wire [13:0] v460; shift_adder #(8, 8, 1, 1, 14, -5, 0) op_460 (v86[7:0], v107[7:0], v460[13:0]); // 1.0
    wire [9:0] v461; shift_adder #(8, 8, 1, 1, 10, 1, 0) op_461 (v119[7:0], v126[7:0], v461[9:0]); // 1.0
    wire [11:0] v462; shift_adder #(8, 8, 1, 1, 12, -3, 0) op_462 (v90[7:0], v90[7:0], v462[11:0]); // 1.0
    wire [9:0] v463; shift_adder #(8, 8, 1, 1, 10, -1, 0) op_463 (v103[7:0], v74[7:0], v463[9:0]); // 1.0
    wire [11:0] v464; shift_adder #(8, 8, 1, 1, 12, -3, 0) op_464 (v115[7:0], v115[7:0], v464[11:0]); // 1.0
    wire [14:0] v465; shift_adder #(8, 8, 1, 1, 15, 6, 1) op_465 (v70[7:0], v112[7:0], v465[14:0]); // 1.0
    wire [9:0] v466; shift_adder #(8, 8, 1, 1, 10, 1, 1) op_466 (v100[7:0], v93[7:0], v466[9:0]); // 1.0
    wire [8:0] v467; shift_adder #(8, 8, 1, 1, 9, 0, 1) op_467 (v111[7:0], v69[7:0], v467[8:0]); // 1.0
    wire [9:0] v468; shift_adder #(8, 8, 1, 1, 10, 1, 1) op_468 (v124[7:0], v109[7:0], v468[9:0]); // 1.0
    wire [9:0] v469; shift_adder #(8, 8, 1, 1, 10, 1, 0) op_469 (v98[7:0], v110[7:0], v469[9:0]); // 1.0
    wire [9:0] v470; shift_adder #(8, 8, 1, 1, 10, -1, 1) op_470 (v66[7:0], v82[7:0], v470[9:0]); // 1.0
    wire [14:0] v471; shift_adder #(8, 8, 1, 1, 15, 6, 0) op_471 (v104[7:0], v81[7:0], v471[14:0]); // 1.0
    wire [13:0] v472; shift_adder #(8, 8, 1, 1, 14, -5, 1) op_472 (v75[7:0], v105[7:0], v472[13:0]); // 1.0
    wire [11:0] v473; shift_adder #(8, 8, 1, 1, 12, -3, 1) op_473 (v90[7:0], v90[7:0], v473[11:0]); // 1.0
    wire [13:0] v474; shift_adder #(8, 8, 1, 1, 14, 5, 1) op_474 (v119[7:0], v68[7:0], v474[13:0]); // 1.0
    wire [11:0] v475; shift_adder #(8, 8, 1, 1, 12, -3, 1) op_475 (v74[7:0], v74[7:0], v475[11:0]); // 1.0
    wire [12:0] v476; shift_adder #(8, 8, 1, 1, 13, 4, 1) op_476 (v65[7:0], v102[7:0], v476[12:0]); // 1.0
    wire [8:0] v477; shift_adder #(8, 8, 1, 1, 9, 0, 0) op_477 (v64[7:0], v71[7:0], v477[8:0]); // 1.0
    wire [10:0] v478; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_478 (v98[7:0], v113[7:0], v478[10:0]); // 1.0
    wire [8:0] v479; shift_adder #(8, 8, 1, 1, 9, 0, 0) op_479 (v88[7:0], v92[7:0], v479[8:0]); // 1.0
    wire [26:0] v480; shift_adder #(8, 8, 1, 1, 27, -18, 1) op_480 (v111[7:0], v111[7:0], v480[26:0]); // 1.0
    wire [13:0] v481; shift_adder #(8, 8, 1, 1, 14, 5, 0) op_481 (v65[7:0], v124[7:0], v481[13:0]); // 1.0
    wire [14:0] v482; shift_adder #(8, 8, 1, 1, 15, 6, 1) op_482 (v79[7:0], v108[7:0], v482[14:0]); // 1.0
    wire [13:0] v483; shift_adder #(8, 8, 1, 1, 14, 5, 0) op_483 (v93[7:0], v72[7:0], v483[13:0]); // 1.0
    wire [19:0] v484; shift_adder #(8, 8, 1, 1, 20, -11, 0) op_484 (v99[7:0], v101[7:0], v484[19:0]); // 1.0
    wire [18:0] v485; shift_adder #(8, 8, 1, 1, 19, -10, 0) op_485 (v118[7:0], v108[7:0], v485[18:0]); // 1.0
    wire [8:0] v486; shift_adder #(8, 8, 1, 1, 9, 0, 1) op_486 (v70[7:0], v93[7:0], v486[8:0]); // 1.0
    wire [10:0] v487; shift_adder #(8, 8, 1, 1, 11, 2, 1) op_487 (v79[7:0], v110[7:0], v487[10:0]); // 1.0
    wire [13:0] v488; shift_adder #(8, 8, 1, 1, 14, -5, 1) op_488 (v89[7:0], v94[7:0], v488[13:0]); // 1.0
    wire [9:0] v489; shift_adder #(8, 8, 1, 1, 10, 1, 1) op_489 (v119[7:0], v88[7:0], v489[9:0]); // 1.0
    wire [8:0] v490; shift_adder #(8, 8, 1, 1, 9, 0, 0) op_490 (v124[7:0], v118[7:0], v490[8:0]); // 1.0
    wire [10:0] v491; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_491 (v78[7:0], v110[7:0], v491[10:0]); // 1.0
    wire [12:0] v492; shift_adder #(8, 8, 1, 1, 13, 4, 1) op_492 (v66[7:0], v90[7:0], v492[12:0]); // 1.0
    wire [17:0] v493; shift_adder #(8, 8, 1, 1, 18, -9, 0) op_493 (v91[7:0], v102[7:0], v493[17:0]); // 1.0
    wire [17:0] v494; shift_adder #(8, 8, 1, 1, 18, -9, 0) op_494 (v127[7:0], v102[7:0], v494[17:0]); // 1.0
    wire [11:0] v495; shift_adder #(8, 8, 1, 1, 12, -3, 0) op_495 (v110[7:0], v110[7:0], v495[11:0]); // 1.0
    wire [12:0] v496; shift_adder #(8, 8, 1, 1, 13, -4, 1) op_496 (v73[7:0], v77[7:0], v496[12:0]); // 1.0
    wire [10:0] v497; shift_adder #(8, 8, 1, 1, 11, 2, 1) op_497 (v87[7:0], v95[7:0], v497[10:0]); // 1.0
    wire [20:0] v498; shift_adder #(8, 8, 1, 1, 21, 12, 0) op_498 (v80[7:0], v80[7:0], v498[20:0]); // 1.0
    wire [13:0] v499; shift_adder #(8, 8, 1, 1, 14, 5, 0) op_499 (v111[7:0], v120[7:0], v499[13:0]); // 1.0
    wire [11:0] v500; shift_adder #(8, 8, 1, 1, 12, -3, 0) op_500 (v127[7:0], v68[7:0], v500[11:0]); // 1.0
    wire [9:0] v501; shift_adder #(8, 8, 1, 1, 10, 1, 0) op_501 (v121[7:0], v107[7:0], v501[9:0]); // 1.0
    wire [11:0] v502; shift_adder #(8, 8, 1, 1, 12, -3, 0) op_502 (v88[7:0], v88[7:0], v502[11:0]); // 1.0
    wire [8:0] v503; shift_adder #(8, 8, 1, 1, 9, 0, 1) op_503 (v68[7:0], v108[7:0], v503[8:0]); // 1.0
    wire [15:0] v504; shift_adder #(8, 8, 1, 1, 16, 7, 1) op_504 (v104[7:0], v86[7:0], v504[15:0]); // 1.0
    wire [10:0] v505; shift_adder #(8, 8, 1, 1, 11, 2, 0) op_505 (v103[7:0], v78[7:0], v505[10:0]); // 1.0
    wire [12:0] v506; shift_adder #(8, 8, 1, 1, 13, -4, 1) op_506 (v121[7:0], v72[7:0], v506[12:0]); // 1.0
    wire [11:0] v507; shift_adder #(8, 8, 1, 1, 12, -3, 1) op_507 (v70[7:0], v70[7:0], v507[11:0]); // 1.0
    wire [8:0] v508; shift_adder #(8, 8, 1, 1, 9, 0, 0) op_508 (v105[7:0], v89[7:0], v508[8:0]); // 1.0
    wire [9:0] v509; shift_adder #(8, 8, 1, 1, 10, -1, 1) op_509 (v127[7:0], v80[7:0], v509[9:0]); // 1.0
    wire [9:0] v510; shift_adder #(8, 8, 1, 1, 10, 1, 0) op_510 (v106[7:0], v113[7:0], v510[9:0]); // 1.0
    wire [34:0] v511; shift_adder #(8, 8, 1, 1, 35, -26, 1) op_511 (v76[7:0], v70[7:0], v511[34:0]); // 1.0
    wire [11:0] v512; shift_adder #(8, 8, 1, 1, 12, 3, 1) op_512 (v116[7:0], v107[7:0], v512[11:0]); // 1.0
    wire [13:0] v513; shift_adder #(8, 8, 1, 1, 14, -5, 0) op_513 (v94[7:0], v64[7:0], v513[13:0]); // 1.0
    wire [13:0] v514; shift_adder #(8, 8, 1, 1, 14, 5, 1) op_514 (v73[7:0], v117[7:0], v514[13:0]); // 1.0
    wire [19:0] v515; shift_adder #(8, 8, 1, 1, 20, -11, 0) op_515 (v87[7:0], v92[7:0], v515[19:0]); // 1.0
    wire [9:0] v516; shift_adder #(8, 8, 1, 1, 10, 1, 0) op_516 (v75[7:0], v73[7:0], v516[9:0]); // 1.0
    wire [25:0] v517; shift_adder #(8, 8, 1, 1, 26, 17, 0) op_517 (v76[7:0], v70[7:0], v517[25:0]); // 1.0
    wire [10:0] v518; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_518 (v85[7:0], v85[7:0], v518[10:0]); // 1.0
    wire [15:0] v519; shift_adder #(8, 8, 1, 1, 16, 7, 1) op_519 (v121[7:0], v64[7:0], v519[15:0]); // 1.0
    wire [9:0] v520; shift_adder #(8, 8, 1, 1, 10, 1, 1) op_520 (v100[7:0], v72[7:0], v520[9:0]); // 1.0
    wire [11:0] v521; shift_adder #(8, 8, 1, 1, 12, -3, 0) op_521 (v87[7:0], v81[7:0], v521[11:0]); // 1.0
    wire [8:0] v522; shift_adder #(8, 8, 1, 1, 9, 0, 0) op_522 (v95[7:0], v102[7:0], v522[8:0]); // 1.0
    wire [11:0] v523; shift_adder #(8, 8, 1, 1, 12, -3, 1) op_523 (v78[7:0], v117[7:0], v523[11:0]); // 1.0
    wire [12:0] v524; shift_adder #(8, 8, 1, 1, 13, -4, 1) op_524 (v65[7:0], v73[7:0], v524[12:0]); // 1.0
    wire [25:0] v525; shift_adder #(8, 8, 1, 1, 26, 17, 0) op_525 (v114[7:0], v64[7:0], v525[25:0]); // 1.0
    wire [14:0] v526; shift_adder #(8, 8, 1, 1, 15, 6, 0) op_526 (v104[7:0], v101[7:0], v526[14:0]); // 1.0
    wire [9:0] v527; shift_adder #(8, 8, 1, 1, 10, -1, 0) op_527 (v104[7:0], v84[7:0], v527[9:0]); // 1.0
    wire [14:0] v528; shift_adder #(8, 8, 1, 1, 15, 6, 0) op_528 (v122[7:0], v77[7:0], v528[14:0]); // 1.0
    wire [23:0] v529; shift_adder #(8, 8, 1, 1, 24, -15, 0) op_529 (v102[7:0], v66[7:0], v529[23:0]); // 1.0
    wire [25:0] v530; shift_adder #(8, 8, 1, 1, 26, 17, 1) op_530 (v109[7:0], v76[7:0], v530[25:0]); // 1.0
    wire [8:0] v531; shift_adder #(8, 8, 1, 1, 9, 0, 1) op_531 (v111[7:0], v122[7:0], v531[8:0]); // 1.0
    wire [11:0] v532; shift_adder #(8, 8, 1, 1, 12, -3, 1) op_532 (v119[7:0], v114[7:0], v532[11:0]); // 1.0
    wire [16:0] v533; shift_adder #(8, 8, 1, 1, 17, 8, 1) op_533 (v109[7:0], v74[7:0], v533[16:0]); // 1.0
    wire [12:0] v534; shift_adder #(8, 8, 1, 1, 13, -4, 0) op_534 (v75[7:0], v66[7:0], v534[12:0]); // 1.0
    wire [17:0] v535; shift_adder #(8, 8, 1, 1, 18, 9, 1) op_535 (v75[7:0], v106[7:0], v535[17:0]); // 1.0
    wire [18:0] v536; shift_adder #(8, 8, 1, 1, 19, -10, 0) op_536 (v127[7:0], v116[7:0], v536[18:0]); // 1.0
    wire [24:0] v537; shift_adder #(8, 8, 1, 1, 25, -16, 0) op_537 (v105[7:0], v116[7:0], v537[24:0]); // 1.0
    wire [8:0] v538; shift_adder #(8, 8, 1, 1, 9, 0, 1) op_538 (v123[7:0], v126[7:0], v538[8:0]); // 1.0
    wire [18:0] v539; shift_adder #(8, 8, 1, 1, 19, -10, 1) op_539 (v118[7:0], v117[7:0], v539[18:0]); // 1.0
    wire [11:0] v540; shift_adder #(8, 8, 1, 1, 12, -3, 1) op_540 (v83[7:0], v83[7:0], v540[11:0]); // 1.0
    wire [11:0] v541; shift_adder #(8, 8, 1, 1, 12, 3, 1) op_541 (v123[7:0], v119[7:0], v541[11:0]); // 1.0
    wire [9:0] v542; shift_adder #(8, 8, 1, 1, 10, -1, 1) op_542 (v122[7:0], v85[7:0], v542[9:0]); // 1.0
    wire [11:0] v543; shift_adder #(8, 8, 1, 1, 12, 3, 0) op_543 (v67[7:0], v89[7:0], v543[11:0]); // 1.0
    wire [11:0] v544; shift_adder #(8, 8, 1, 1, 12, 3, 0) op_544 (v106[7:0], v98[7:0], v544[11:0]); // 1.0
    wire [16:0] v545; shift_adder #(8, 8, 1, 1, 17, -8, 1) op_545 (v94[7:0], v90[7:0], v545[16:0]); // 1.0
    wire [15:0] v546; shift_adder #(8, 8, 1, 1, 16, -7, 1) op_546 (v121[7:0], v67[7:0], v546[15:0]); // 1.0
    wire [18:0] v547; shift_adder #(8, 8, 1, 1, 19, 10, 0) op_547 (v84[7:0], v115[7:0], v547[18:0]); // 1.0
    wire [9:0] v548; shift_adder #(8, 8, 1, 1, 10, -1, 0) op_548 (v115[7:0], v90[7:0], v548[9:0]); // 1.0
    wire [9:0] v549; shift_adder #(8, 8, 1, 1, 10, 1, 1) op_549 (v70[7:0], v93[7:0], v549[9:0]); // 1.0
    wire [11:0] v550; shift_adder #(8, 8, 1, 1, 12, -3, 1) op_550 (v76[7:0], v76[7:0], v550[11:0]); // 1.0
    wire [16:0] v551; shift_adder #(8, 8, 1, 1, 17, -8, 0) op_551 (v91[7:0], v85[7:0], v551[16:0]); // 1.0
    wire [11:0] v552; shift_adder #(8, 8, 1, 1, 12, 3, 0) op_552 (v102[7:0], v67[7:0], v552[11:0]); // 1.0
    wire [11:0] v553; shift_adder #(8, 8, 1, 1, 12, -3, 1) op_553 (v100[7:0], v100[7:0], v553[11:0]); // 1.0
    wire [9:0] v554; shift_adder #(8, 8, 1, 1, 10, -1, 0) op_554 (v65[7:0], v80[7:0], v554[9:0]); // 1.0
    wire [13:0] v555; shift_adder #(8, 8, 1, 1, 14, -5, 0) op_555 (v122[7:0], v85[7:0], v555[13:0]); // 1.0
    wire [8:0] v556; shift_adder #(8, 8, 1, 1, 9, 0, 0) op_556 (v93[7:0], v71[7:0], v556[8:0]); // 1.0
    wire [14:0] v557; shift_adder #(8, 8, 1, 1, 15, -6, 0) op_557 (v113[7:0], v68[7:0], v557[14:0]); // 1.0
    wire [18:0] v558; shift_adder #(8, 8, 1, 1, 19, -10, 1) op_558 (v65[7:0], v82[7:0], v558[18:0]); // 1.0
    wire [23:0] v559; shift_adder #(8, 8, 1, 1, 24, -15, 1) op_559 (v104[7:0], v115[7:0], v559[23:0]); // 1.0
    wire [19:0] v560; shift_adder #(8, 8, 1, 1, 20, 11, 0) op_560 (v92[7:0], v121[7:0], v560[19:0]); // 1.0
    wire [8:0] v561; shift_adder #(8, 8, 1, 1, 9, 0, 0) op_561 (v96[7:0], v79[7:0], v561[8:0]); // 1.0
    wire [17:0] v562; shift_adder #(8, 8, 1, 1, 18, -9, 0) op_562 (v87[7:0], v67[7:0], v562[17:0]); // 1.0
    wire [10:0] v563; shift_adder #(8, 8, 1, 1, 11, 2, 0) op_563 (v114[7:0], v84[7:0], v563[10:0]); // 1.0
    wire [22:0] v564; shift_adder #(8, 8, 1, 1, 23, -14, 1) op_564 (v98[7:0], v98[7:0], v564[22:0]); // 1.0
    wire [9:0] v565; shift_adder #(8, 8, 1, 1, 10, 1, 0) op_565 (v97[7:0], v73[7:0], v565[9:0]); // 1.0
    wire [15:0] v566; shift_adder #(8, 8, 1, 1, 16, 7, 0) op_566 (v96[7:0], v117[7:0], v566[15:0]); // 1.0
    wire [9:0] v567; shift_adder #(8, 8, 1, 1, 10, -1, 0) op_567 (v107[7:0], v64[7:0], v567[9:0]); // 1.0
    wire [8:0] v568; shift_adder #(8, 8, 1, 1, 9, 0, 1) op_568 (v70[7:0], v98[7:0], v568[8:0]); // 1.0
    wire [9:0] v569; shift_adder #(8, 8, 1, 1, 10, 1, 0) op_569 (v103[7:0], v73[7:0], v569[9:0]); // 1.0
    wire [10:0] v570; shift_adder #(8, 8, 1, 1, 11, 2, 0) op_570 (v107[7:0], v124[7:0], v570[10:0]); // 1.0
    wire [13:0] v571; shift_adder #(8, 8, 1, 1, 14, -5, 0) op_571 (v85[7:0], v71[7:0], v571[13:0]); // 1.0
    wire [9:0] v572; shift_adder #(8, 8, 1, 1, 10, 1, 0) op_572 (v94[7:0], v114[7:0], v572[9:0]); // 1.0
    wire [12:0] v573; shift_adder #(8, 8, 1, 1, 13, 4, 0) op_573 (v109[7:0], v80[7:0], v573[12:0]); // 1.0
    wire [10:0] v574; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_574 (v112[7:0], v76[7:0], v574[10:0]); // 1.0
    wire [8:0] v575; shift_adder #(8, 8, 1, 1, 9, 0, 1) op_575 (v105[7:0], v86[7:0], v575[8:0]); // 1.0
    wire [9:0] v576; shift_adder #(8, 8, 1, 1, 10, 1, 0) op_576 (v114[7:0], v84[7:0], v576[9:0]); // 1.0
    wire [10:0] v577; shift_adder #(8, 8, 1, 1, 11, -2, 1) op_577 (v101[7:0], v71[7:0], v577[10:0]); // 1.0
    wire [12:0] v578; shift_adder #(8, 8, 1, 1, 13, -4, 1) op_578 (v83[7:0], v72[7:0], v578[12:0]); // 1.0
    wire [11:0] v579; shift_adder #(8, 8, 1, 1, 12, -3, 0) op_579 (v118[7:0], v118[7:0], v579[11:0]); // 1.0
    wire [22:0] v580; shift_adder #(8, 8, 1, 1, 23, 14, 0) op_580 (v126[7:0], v80[7:0], v580[22:0]); // 1.0
    wire [10:0] v581; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_581 (v125[7:0], v86[7:0], v581[10:0]); // 1.0
    wire [11:0] v582; shift_adder #(8, 8, 1, 1, 12, -3, 1) op_582 (v114[7:0], v107[7:0], v582[11:0]); // 1.0
    wire [15:0] v583; shift_adder #(8, 8, 1, 1, 16, -7, 0) op_583 (v65[7:0], v85[7:0], v583[15:0]); // 1.0
    wire [9:0] v584; shift_adder #(8, 8, 1, 1, 10, 1, 1) op_584 (v118[7:0], v71[7:0], v584[9:0]); // 1.0
    wire [9:0] v585; shift_adder #(8, 8, 1, 1, 10, -1, 1) op_585 (v83[7:0], v120[7:0], v585[9:0]); // 1.0
    wire [11:0] v586; shift_adder #(8, 8, 1, 1, 12, -3, 1) op_586 (v75[7:0], v106[7:0], v586[11:0]); // 1.0
    wire [21:0] v587; shift_adder #(8, 8, 1, 1, 22, 13, 0) op_587 (v110[7:0], v90[7:0], v587[21:0]); // 1.0
    wire [33:0] v588; shift_adder #(8, 8, 1, 1, 34, 25, 0) op_588 (v80[7:0], v87[7:0], v588[33:0]); // 1.0
    wire [11:0] v589; shift_adder #(8, 8, 1, 1, 12, -3, 0) op_589 (v89[7:0], v68[7:0], v589[11:0]); // 1.0
    wire [13:0] v590; shift_adder #(8, 8, 1, 1, 14, -5, 1) op_590 (v95[7:0], v89[7:0], v590[13:0]); // 1.0
    wire [31:0] v591; shift_adder #(8, 8, 1, 1, 32, -23, 1) op_591 (v67[7:0], v106[7:0], v591[31:0]); // 1.0
    wire [9:0] v592; shift_adder #(8, 8, 1, 1, 10, 1, 1) op_592 (v93[7:0], v108[7:0], v592[9:0]); // 1.0
    wire [27:0] v593; shift_adder #(8, 8, 1, 1, 28, 19, 1) op_593 (v91[7:0], v77[7:0], v593[27:0]); // 1.0
    wire [15:0] v594; shift_adder #(8, 8, 1, 1, 16, -7, 0) op_594 (v117[7:0], v117[7:0], v594[15:0]); // 1.0
    wire [24:0] v595; shift_adder #(8, 8, 1, 1, 25, 16, 0) op_595 (v112[7:0], v115[7:0], v595[24:0]); // 1.0
    wire [15:0] v596; shift_adder #(8, 8, 1, 1, 16, -7, 0) op_596 (v125[7:0], v87[7:0], v596[15:0]); // 1.0
    wire [18:0] v597; shift_adder #(8, 8, 1, 1, 19, -10, 1) op_597 (v127[7:0], v102[7:0], v597[18:0]); // 1.0
    wire [12:0] v598; shift_adder #(8, 8, 1, 1, 13, -4, 1) op_598 (v67[7:0], v113[7:0], v598[12:0]); // 1.0
    wire [20:0] v599; shift_adder #(8, 8, 1, 1, 21, -12, 0) op_599 (v97[7:0], v91[7:0], v599[20:0]); // 1.0
    wire [10:0] v600; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_600 (v125[7:0], v92[7:0], v600[10:0]); // 1.0
    wire [12:0] v601; shift_adder #(8, 8, 1, 1, 13, 4, 0) op_601 (v114[7:0], v125[7:0], v601[12:0]); // 1.0
    wire [10:0] v602; shift_adder #(8, 8, 1, 1, 11, 2, 0) op_602 (v66[7:0], v74[7:0], v602[10:0]); // 1.0
    wire [13:0] v603; shift_adder #(8, 8, 1, 1, 14, -5, 1) op_603 (v121[7:0], v72[7:0], v603[13:0]); // 1.0
    wire [19:0] v604; shift_adder #(8, 8, 1, 1, 20, 11, 0) op_604 (v112[7:0], v96[7:0], v604[19:0]); // 1.0
    wire [29:0] v605; shift_adder #(8, 8, 1, 1, 30, 21, 1) op_605 (v106[7:0], v122[7:0], v605[29:0]); // 1.0
    wire [9:0] v606; shift_adder #(8, 8, 1, 1, 10, -1, 1) op_606 (v113[7:0], v76[7:0], v606[9:0]); // 1.0
    wire [10:0] v607; shift_adder #(8, 8, 1, 1, 11, 2, 0) op_607 (v124[7:0], v69[7:0], v607[10:0]); // 1.0
    wire [32:0] v608; shift_adder #(8, 8, 1, 1, 33, -24, 1) op_608 (v124[7:0], v89[7:0], v608[32:0]); // 1.0
    wire [9:0] v609; shift_adder #(8, 8, 1, 1, 10, -1, 1) op_609 (v104[7:0], v93[7:0], v609[9:0]); // 1.0
    wire [9:0] v610; shift_adder #(8, 8, 1, 1, 10, -1, 1) op_610 (v120[7:0], v77[7:0], v610[9:0]); // 1.0
    wire [24:0] v611; shift_adder #(8, 8, 1, 1, 25, -16, 1) op_611 (v85[7:0], v89[7:0], v611[24:0]); // 1.0
    wire [10:0] v612; shift_adder #(8, 8, 1, 1, 11, 2, 0) op_612 (v67[7:0], v105[7:0], v612[10:0]); // 1.0
    wire [26:0] v613; shift_adder #(8, 8, 1, 1, 27, -18, 0) op_613 (v112[7:0], v78[7:0], v613[26:0]); // 1.0
    wire [11:0] v614; shift_adder #(8, 8, 1, 1, 12, -3, 1) op_614 (v101[7:0], v101[7:0], v614[11:0]); // 1.0
    wire [16:0] v615; shift_adder #(8, 8, 1, 1, 17, -8, 0) op_615 (v119[7:0], v73[7:0], v615[16:0]); // 1.0
    wire [10:0] v616; shift_adder #(8, 8, 1, 1, 11, 2, 0) op_616 (v73[7:0], v81[7:0], v616[10:0]); // 1.0
    wire [21:0] v617; shift_adder #(8, 8, 1, 1, 22, 13, 0) op_617 (v103[7:0], v110[7:0], v617[21:0]); // 1.0
    wire [27:0] v618; shift_adder #(8, 8, 1, 1, 28, 19, 0) op_618 (v121[7:0], v91[7:0], v618[27:0]); // 1.0
    wire [18:0] v619; shift_adder #(8, 8, 1, 1, 19, -10, 1) op_619 (v71[7:0], v64[7:0], v619[18:0]); // 1.0
    wire [8:0] v620; shift_adder #(8, 8, 1, 1, 9, 0, 1) op_620 (v97[7:0], v73[7:0], v620[8:0]); // 1.0
    wire [8:0] v621; shift_adder #(8, 8, 1, 1, 9, 0, 0) op_621 (v99[7:0], v72[7:0], v621[8:0]); // 1.0
    wire [10:0] v622; shift_adder #(8, 8, 1, 1, 11, 2, 0) op_622 (v105[7:0], v77[7:0], v622[10:0]); // 1.0
    wire [21:0] v623; shift_adder #(8, 8, 1, 1, 22, -13, 0) op_623 (v123[7:0], v106[7:0], v623[21:0]); // 1.0
    wire [20:0] v624; shift_adder #(8, 8, 1, 1, 21, 12, 0) op_624 (v118[7:0], v113[7:0], v624[20:0]); // 1.0
    wire [12:0] v625; shift_adder #(8, 8, 1, 1, 13, -4, 1) op_625 (v83[7:0], v102[7:0], v625[12:0]); // 1.0
    wire [9:0] v626; shift_adder #(8, 8, 1, 1, 10, 1, 0) op_626 (v67[7:0], v94[7:0], v626[9:0]); // 1.0
    wire [8:0] v627; shift_adder #(8, 8, 1, 1, 9, 0, 1) op_627 (v109[7:0], v73[7:0], v627[8:0]); // 1.0
    wire [19:0] v628; shift_adder #(8, 8, 1, 1, 20, 11, 0) op_628 (v90[7:0], v125[7:0], v628[19:0]); // 1.0
    wire [11:0] v629; shift_adder #(8, 8, 1, 1, 12, 3, 0) op_629 (v121[7:0], v117[7:0], v629[11:0]); // 1.0
    wire [14:0] v630; shift_adder #(8, 8, 1, 1, 15, -6, 1) op_630 (v116[7:0], v120[7:0], v630[14:0]); // 1.0
    wire [12:0] v631; shift_adder #(8, 8, 1, 1, 13, 4, 0) op_631 (v98[7:0], v120[7:0], v631[12:0]); // 1.0
    wire [9:0] v632; shift_adder #(8, 8, 1, 1, 10, 1, 1) op_632 (v114[7:0], v79[7:0], v632[9:0]); // 1.0
    wire [17:0] v633; shift_adder #(8, 8, 1, 1, 18, 9, 0) op_633 (v97[7:0], v110[7:0], v633[17:0]); // 1.0
    wire [15:0] v634; shift_adder #(8, 8, 1, 1, 16, -7, 0) op_634 (v108[7:0], v73[7:0], v634[15:0]); // 1.0
    wire [22:0] v635; shift_adder #(8, 8, 1, 1, 23, 14, 0) op_635 (v114[7:0], v74[7:0], v635[22:0]); // 1.0
    wire [10:0] v636; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_636 (v85[7:0], v103[7:0], v636[10:0]); // 1.0
    wire [8:0] v637; shift_adder #(8, 8, 1, 1, 9, 0, 0) op_637 (v79[7:0], v71[7:0], v637[8:0]); // 1.0
    wire [13:0] v638; shift_adder #(8, 8, 1, 1, 14, -5, 0) op_638 (v93[7:0], v115[7:0], v638[13:0]); // 1.0
    wire [9:0] v639; shift_adder #(8, 8, 1, 1, 10, -1, 0) op_639 (v74[7:0], v64[7:0], v639[9:0]); // 1.0
    wire [18:0] v640; shift_adder #(8, 8, 1, 1, 19, 10, 1) op_640 (v79[7:0], v86[7:0], v640[18:0]); // 1.0
    wire [30:0] v641; shift_adder #(8, 8, 1, 1, 31, 22, 1) op_641 (v125[7:0], v92[7:0], v641[30:0]); // 1.0
    wire [11:0] v642; shift_adder #(8, 8, 1, 1, 12, -3, 0) op_642 (v84[7:0], v76[7:0], v642[11:0]); // 1.0
    wire [9:0] v643; shift_adder #(8, 8, 1, 1, 10, -1, 1) op_643 (v106[7:0], v81[7:0], v643[9:0]); // 1.0
    wire [10:0] v644; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_644 (v88[7:0], v115[7:0], v644[10:0]); // 1.0
    wire [12:0] v645; shift_adder #(8, 8, 1, 1, 13, -4, 0) op_645 (v68[7:0], v68[7:0], v645[12:0]); // 1.0
    wire [12:0] v646; shift_adder #(8, 8, 1, 1, 13, 4, 0) op_646 (v72[7:0], v121[7:0], v646[12:0]); // 1.0
    wire [9:0] v647; shift_adder #(8, 8, 1, 1, 10, 1, 0) op_647 (v116[7:0], v92[7:0], v647[9:0]); // 1.0
    wire [9:0] v648; shift_adder #(8, 8, 1, 1, 10, -1, 0) op_648 (v86[7:0], v67[7:0], v648[9:0]); // 1.0
    wire [14:0] v649; shift_adder #(8, 8, 1, 1, 15, -6, 1) op_649 (v84[7:0], v86[7:0], v649[14:0]); // 1.0
    wire [11:0] v650; shift_adder #(8, 8, 1, 1, 12, -3, 0) op_650 (v119[7:0], v92[7:0], v650[11:0]); // 1.0
    wire [8:0] v651; shift_adder #(8, 8, 1, 1, 9, 0, 0) op_651 (v93[7:0], v75[7:0], v651[8:0]); // 1.0
    wire [14:0] v652; shift_adder #(8, 8, 1, 1, 15, -6, 0) op_652 (v122[7:0], v113[7:0], v652[14:0]); // 1.0
    wire [10:0] v653; shift_adder #(8, 8, 1, 1, 11, 2, 0) op_653 (v98[7:0], v122[7:0], v653[10:0]); // 1.0
    wire [12:0] v654; shift_adder #(8, 8, 1, 1, 13, -4, 1) op_654 (v116[7:0], v116[7:0], v654[12:0]); // 1.0
    wire [15:0] v655; shift_adder #(8, 8, 1, 1, 16, -7, 0) op_655 (v65[7:0], v94[7:0], v655[15:0]); // 1.0
    wire [21:0] v656; shift_adder #(8, 8, 1, 1, 22, -13, 0) op_656 (v69[7:0], v69[7:0], v656[21:0]); // 1.0
    wire [11:0] v657; shift_adder #(8, 8, 1, 1, 12, -3, 0) op_657 (v87[7:0], v121[7:0], v657[11:0]); // 1.0
    wire [13:0] v658; shift_adder #(8, 8, 1, 1, 14, -5, 0) op_658 (v71[7:0], v108[7:0], v658[13:0]); // 1.0
    wire [10:0] v659; shift_adder #(8, 8, 1, 1, 11, -2, 1) op_659 (v124[7:0], v92[7:0], v659[10:0]); // 1.0
    wire [12:0] v660; shift_adder #(8, 8, 1, 1, 13, -4, 0) op_660 (v82[7:0], v90[7:0], v660[12:0]); // 1.0
    wire [10:0] v661; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_661 (v103[7:0], v106[7:0], v661[10:0]); // 1.0
    wire [10:0] v662; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_662 (v106[7:0], v98[7:0], v662[10:0]); // 1.0
    wire [8:0] v663; shift_adder #(8, 8, 1, 1, 9, 0, 0) op_663 (v112[7:0], v110[7:0], v663[8:0]); // 1.0
    wire [11:0] v664; shift_adder #(8, 8, 1, 1, 12, 3, 0) op_664 (v93[7:0], v101[7:0], v664[11:0]); // 1.0
    wire [13:0] v665; shift_adder #(8, 8, 1, 1, 14, 5, 0) op_665 (v77[7:0], v81[7:0], v665[13:0]); // 1.0
    wire [9:0] v666; shift_adder #(8, 8, 1, 1, 10, 1, 0) op_666 (v66[7:0], v99[7:0], v666[9:0]); // 1.0
    wire [16:0] v667; shift_adder #(8, 8, 1, 1, 17, -8, 0) op_667 (v95[7:0], v80[7:0], v667[16:0]); // 1.0
    wire [11:0] v668; shift_adder #(8, 8, 1, 1, 12, 3, 0) op_668 (v92[7:0], v81[7:0], v668[11:0]); // 1.0
    wire [9:0] v669; shift_adder #(8, 8, 1, 1, 10, 1, 0) op_669 (v112[7:0], v127[7:0], v669[9:0]); // 1.0
    wire [34:0] v670; shift_adder #(8, 8, 1, 1, 35, -26, 1) op_670 (v82[7:0], v70[7:0], v670[34:0]); // 1.0
    wire [10:0] v671; shift_adder #(8, 8, 1, 1, 11, 2, 0) op_671 (v106[7:0], v90[7:0], v671[10:0]); // 1.0
    wire [10:0] v672; shift_adder #(8, 8, 1, 1, 11, 2, 0) op_672 (v122[7:0], v67[7:0], v672[10:0]); // 1.0
    wire [12:0] v673; shift_adder #(8, 8, 1, 1, 13, 4, 0) op_673 (v112[7:0], v77[7:0], v673[12:0]); // 1.0
    wire [14:0] v674; shift_adder #(8, 8, 1, 1, 15, 6, 0) op_674 (v104[7:0], v119[7:0], v674[14:0]); // 1.0
    wire [10:0] v675; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_675 (v96[7:0], v113[7:0], v675[10:0]); // 1.0
    wire [10:0] v676; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_676 (v124[7:0], v117[7:0], v676[10:0]); // 1.0
    wire [16:0] v677; shift_adder #(8, 8, 1, 1, 17, -8, 1) op_677 (v96[7:0], v67[7:0], v677[16:0]); // 1.0
    wire [9:0] v678; shift_adder #(8, 8, 1, 1, 10, 1, 0) op_678 (v99[7:0], v77[7:0], v678[9:0]); // 1.0
    wire [10:0] v679; shift_adder #(8, 8, 1, 1, 11, 2, 0) op_679 (v89[7:0], v74[7:0], v679[10:0]); // 1.0
    wire [23:0] v680; shift_adder #(8, 8, 1, 1, 24, -15, 0) op_680 (v75[7:0], v80[7:0], v680[23:0]); // 1.0
    wire [17:0] v681; shift_adder #(8, 8, 1, 1, 18, -9, 0) op_681 (v106[7:0], v90[7:0], v681[17:0]); // 1.0
    wire [17:0] v682; shift_adder #(8, 8, 1, 1, 18, 9, 1) op_682 (v96[7:0], v104[7:0], v682[17:0]); // 1.0
    wire [34:0] v683; shift_adder #(8, 8, 1, 1, 35, -26, 1) op_683 (v113[7:0], v99[7:0], v683[34:0]); // 1.0
    wire [31:0] v684; shift_adder #(8, 8, 1, 1, 32, 23, 0) op_684 (v110[7:0], v80[7:0], v684[31:0]); // 1.0
    wire [10:0] v685; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_685 (v83[7:0], v80[7:0], v685[10:0]); // 1.0
    wire [11:0] v686; shift_adder #(8, 8, 1, 1, 12, -3, 0) op_686 (v80[7:0], v123[7:0], v686[11:0]); // 1.0
    wire [13:0] v687; shift_adder #(8, 8, 1, 1, 14, -5, 0) op_687 (v124[7:0], v115[7:0], v687[13:0]); // 1.0
    wire [10:0] v688; shift_adder #(8, 8, 1, 1, 11, -2, 1) op_688 (v122[7:0], v102[7:0], v688[10:0]); // 1.0
    wire [16:0] v689; shift_adder #(8, 8, 1, 1, 17, 8, 1) op_689 (v99[7:0], v94[7:0], v689[16:0]); // 1.0
    wire [14:0] v690; shift_adder #(8, 8, 1, 1, 15, 6, 0) op_690 (v101[7:0], v116[7:0], v690[14:0]); // 1.0
    wire [11:0] v691; shift_adder #(8, 8, 1, 1, 12, 3, 0) op_691 (v98[7:0], v72[7:0], v691[11:0]); // 1.0
    wire [10:0] v692; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_692 (v120[7:0], v66[7:0], v692[10:0]); // 1.0
    wire [8:0] v693; shift_adder #(8, 8, 1, 1, 9, 0, 0) op_693 (v107[7:0], v81[7:0], v693[8:0]); // 1.0
    wire [10:0] v694; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_694 (v89[7:0], v127[7:0], v694[10:0]); // 1.0
    wire [14:0] v695; shift_adder #(8, 8, 1, 1, 15, -6, 0) op_695 (v121[7:0], v76[7:0], v695[14:0]); // 1.0
    wire [10:0] v696; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_696 (v67[7:0], v71[7:0], v696[10:0]); // 1.0
    wire [14:0] v697; shift_adder #(8, 8, 1, 1, 15, 6, 0) op_697 (v110[7:0], v75[7:0], v697[14:0]); // 1.0
    wire [13:0] v698; shift_adder #(8, 8, 1, 1, 14, 5, 0) op_698 (v113[7:0], v98[7:0], v698[13:0]); // 1.0
    wire [9:0] v699; shift_adder #(8, 8, 1, 1, 10, -1, 0) op_699 (v112[7:0], v71[7:0], v699[9:0]); // 1.0
    wire [14:0] v700; shift_adder #(8, 8, 1, 1, 15, -6, 0) op_700 (v120[7:0], v79[7:0], v700[14:0]); // 1.0
    wire [10:0] v701; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_701 (v118[7:0], v124[7:0], v701[10:0]); // 1.0
    wire [10:0] v702; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_702 (v82[7:0], v86[7:0], v702[10:0]); // 1.0
    wire [14:0] v703; shift_adder #(8, 8, 1, 1, 15, -6, 0) op_703 (v95[7:0], v70[7:0], v703[14:0]); // 1.0
    wire [9:0] v704; shift_adder #(8, 8, 1, 1, 10, -1, 0) op_704 (v78[7:0], v81[7:0], v704[9:0]); // 1.0
    wire [9:0] v705; shift_adder #(8, 8, 1, 1, 10, 1, 0) op_705 (v88[7:0], v72[7:0], v705[9:0]); // 1.0
    wire [14:0] v706; shift_adder #(8, 8, 1, 1, 15, 6, 0) op_706 (v127[7:0], v102[7:0], v706[14:0]); // 1.0
    wire [9:0] v707; shift_adder #(8, 8, 1, 1, 10, 1, 0) op_707 (v86[7:0], v111[7:0], v707[9:0]); // 1.0
    wire [10:0] v708; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_708 (v88[7:0], v77[7:0], v708[10:0]); // 1.0
    wire [11:0] v709; shift_adder #(8, 8, 1, 1, 12, -3, 0) op_709 (v90[7:0], v91[7:0], v709[11:0]); // 1.0
    wire [15:0] v710; shift_adder #(8, 8, 1, 1, 16, -7, 0) op_710 (v93[7:0], v105[7:0], v710[15:0]); // 1.0
    wire [15:0] v711; shift_adder #(8, 8, 1, 1, 16, 7, 0) op_711 (v74[7:0], v98[7:0], v711[15:0]); // 1.0
    wire [10:0] v712; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_712 (v88[7:0], v108[7:0], v712[10:0]); // 1.0
    wire [28:0] v713; shift_adder #(8, 8, 1, 1, 29, -20, 1) op_713 (v85[7:0], v83[7:0], v713[28:0]); // 1.0
    wire [10:0] v714; shift_adder #(8, 8, 1, 1, 11, 2, 0) op_714 (v96[7:0], v90[7:0], v714[10:0]); // 1.0
    wire [12:0] v715; shift_adder #(8, 8, 1, 1, 13, -4, 0) op_715 (v100[7:0], v86[7:0], v715[12:0]); // 1.0
    wire [9:0] v716; shift_adder #(8, 8, 1, 1, 10, 1, 1) op_716 (v78[7:0], v77[7:0], v716[9:0]); // 1.0
    wire [9:0] v717; shift_adder #(8, 8, 1, 1, 10, 1, 0) op_717 (v91[7:0], v104[7:0], v717[9:0]); // 1.0
    wire [12:0] v718; shift_adder #(8, 8, 1, 1, 13, -4, 0) op_718 (v90[7:0], v114[7:0], v718[12:0]); // 1.0
    wire [11:0] v719; shift_adder #(8, 8, 1, 1, 12, 3, 0) op_719 (v84[7:0], v64[7:0], v719[11:0]); // 1.0
    wire [26:0] v720; shift_adder #(8, 8, 1, 1, 27, 18, 0) op_720 (v117[7:0], v122[7:0], v720[26:0]); // 1.0
    wire [10:0] v721; shift_adder #(8, 8, 1, 1, 11, 2, 0) op_721 (v64[7:0], v75[7:0], v721[10:0]); // 1.0
    wire [9:0] v722; shift_adder #(8, 8, 1, 1, 10, 1, 0) op_722 (v79[7:0], v76[7:0], v722[9:0]); // 1.0
    wire [10:0] v723; shift_adder #(8, 8, 1, 1, 11, 2, 0) op_723 (v114[7:0], v111[7:0], v723[10:0]); // 1.0
    wire [8:0] v724; shift_adder #(8, 8, 1, 1, 9, 0, 0) op_724 (v69[7:0], v113[7:0], v724[8:0]); // 1.0
    wire [23:0] v725; shift_adder #(8, 8, 1, 1, 24, -15, 0) op_725 (v80[7:0], v109[7:0], v725[23:0]); // 1.0
    wire [32:0] v726; shift_adder #(8, 8, 1, 1, 33, -24, 1) op_726 (v115[7:0], v117[7:0], v726[32:0]); // 1.0
    wire [9:0] v727; shift_adder #(8, 8, 1, 1, 10, -1, 0) op_727 (v85[7:0], v78[7:0], v727[9:0]); // 1.0
    wire [10:0] v728; shift_adder #(8, 8, 1, 1, 11, 2, 0) op_728 (v79[7:0], v121[7:0], v728[10:0]); // 1.0
    wire [10:0] v729; shift_adder #(8, 8, 1, 1, 11, 2, 0) op_729 (v98[7:0], v126[7:0], v729[10:0]); // 1.0
    wire [9:0] v730; shift_adder #(8, 8, 1, 1, 10, 1, 0) op_730 (v125[7:0], v95[7:0], v730[9:0]); // 1.0
    wire [15:0] v731; shift_adder #(8, 8, 1, 1, 16, -7, 0) op_731 (v69[7:0], v101[7:0], v731[15:0]); // 1.0
    wire [18:0] v732; shift_adder #(8, 8, 1, 1, 19, 10, 0) op_732 (v107[7:0], v83[7:0], v732[18:0]); // 1.0
    wire [14:0] v733; shift_adder #(8, 8, 1, 1, 15, -6, 0) op_733 (v105[7:0], v71[7:0], v733[14:0]); // 1.0
    wire [11:0] v734; shift_adder #(8, 8, 1, 1, 12, 3, 0) op_734 (v87[7:0], v68[7:0], v734[11:0]); // 1.0
    wire [12:0] v735; shift_adder #(8, 8, 1, 1, 13, -4, 0) op_735 (v125[7:0], v74[7:0], v735[12:0]); // 1.0
    wire [10:0] v736; shift_adder #(8, 8, 1, 1, 11, 2, 0) op_736 (v126[7:0], v119[7:0], v736[10:0]); // 1.0
    wire [19:0] v737; shift_adder #(8, 8, 1, 1, 20, 11, 0) op_737 (v76[7:0], v74[7:0], v737[19:0]); // 1.0
    wire [10:0] v738; shift_adder #(8, 8, 1, 1, 11, 2, 0) op_738 (v88[7:0], v98[7:0], v738[10:0]); // 1.0
    wire [9:0] v739; shift_adder #(8, 8, 1, 1, 10, 1, 0) op_739 (v122[7:0], v105[7:0], v739[9:0]); // 1.0
    wire [10:0] v740; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_740 (v121[7:0], v118[7:0], v740[10:0]); // 1.0
    wire [17:0] v741; shift_adder #(8, 8, 1, 1, 18, -9, 0) op_741 (v68[7:0], v84[7:0], v741[17:0]); // 1.0
    wire [12:0] v742; shift_adder #(8, 8, 1, 1, 13, -4, 0) op_742 (v116[7:0], v120[7:0], v742[12:0]); // 1.0
    wire [21:0] v743; shift_adder #(8, 8, 1, 1, 22, 13, 0) op_743 (v67[7:0], v79[7:0], v743[21:0]); // 1.0
    wire [12:0] v744; shift_adder #(8, 8, 1, 1, 13, -4, 0) op_744 (v82[7:0], v76[7:0], v744[12:0]); // 1.0
    wire [10:0] v745; shift_adder #(8, 8, 1, 1, 11, 2, 0) op_745 (v90[7:0], v118[7:0], v745[10:0]); // 1.0
    wire [9:0] v746; shift_adder #(8, 8, 1, 1, 10, -1, 0) op_746 (v65[7:0], v67[7:0], v746[9:0]); // 1.0
    wire [10:0] v747; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_747 (v118[7:0], v101[7:0], v747[10:0]); // 1.0
    wire [9:0] v748; shift_adder #(8, 8, 1, 1, 10, 1, 0) op_748 (v108[7:0], v84[7:0], v748[9:0]); // 1.0
    wire [8:0] v749; shift_adder #(8, 8, 1, 1, 9, 0, 0) op_749 (v89[7:0], v95[7:0], v749[8:0]); // 1.0
    wire [10:0] v750; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_750 (v74[7:0], v108[7:0], v750[10:0]); // 1.0
    wire [16:0] v751; shift_adder #(8, 8, 1, 1, 17, 8, 0) op_751 (v82[7:0], v95[7:0], v751[16:0]); // 1.0
    wire [10:0] v752; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_752 (v98[7:0], v70[7:0], v752[10:0]); // 1.0
    wire [22:0] v753; shift_adder #(8, 8, 1, 1, 23, 14, 0) op_753 (v90[7:0], v68[7:0], v753[22:0]); // 1.0
    wire [8:0] v754; shift_adder #(8, 8, 1, 1, 9, 0, 0) op_754 (v107[7:0], v75[7:0], v754[8:0]); // 1.0
    wire [12:0] v755; shift_adder #(8, 8, 1, 1, 13, -4, 0) op_755 (v68[7:0], v83[7:0], v755[12:0]); // 1.0
    wire [10:0] v756; shift_adder #(8, 8, 1, 1, 11, -2, 0) op_756 (v66[7:0], v123[7:0], v756[10:0]); // 1.0
    wire [16:0] v757; shift_adder #(8, 8, 1, 1, 17, 8, 0) op_757 (v119[7:0], v122[7:0], v757[16:0]); // 1.0
    wire [8:0] v758; shift_adder #(8, 8, 1, 1, 9, 0, 0) op_758 (v86[7:0], v71[7:0], v758[8:0]); // 1.0
    wire [16:0] v759; shift_adder #(8, 8, 1, 1, 17, -8, 0) op_759 (v75[7:0], v103[7:0], v759[16:0]); // 1.0
    wire [20:0] v760; shift_adder #(8, 8, 1, 1, 21, 12, 0) op_760 (v117[7:0], v104[7:0], v760[20:0]); // 1.0
    wire [37:0] v761; shift_adder #(8, 8, 1, 1, 38, -29, 1) op_761 (v97[7:0], v114[7:0], v761[37:0]); // 1.0
    wire [11:0] v762; shift_adder #(8, 8, 1, 1, 12, -3, 0) op_762 (v91[7:0], v116[7:0], v762[11:0]); // 1.0
    wire [9:0] v763; shift_adder #(8, 8, 1, 1, 10, -1, 0) op_763 (v86[7:0], v89[7:0], v763[9:0]); // 1.0
    wire [19:0] v764; shift_adder #(8, 8, 1, 1, 20, -11, 0) op_764 (v82[7:0], v110[7:0], v764[19:0]); // 1.0
    wire [13:0] v765; shift_adder #(8, 8, 1, 1, 14, 5, 0) op_765 (v64[7:0], v92[7:0], v765[13:0]); // 1.0
    wire [22:0] v766; shift_adder #(8, 8, 1, 1, 23, -14, 1) op_766 (v108[7:0], v91[7:0], v766[22:0]); // 1.0
    wire [14:0] v767; shift_adder #(8, 8, 1, 1, 15, 6, 0) op_767 (v81[7:0], v75[7:0], v767[14:0]); // 1.0
    wire [10:0] v768; shift_adder #(8, 8, 1, 1, 11, 2, 0) op_768 (v87[7:0], v115[7:0], v768[10:0]); // 1.0
    wire [10:0] v769; shift_adder #(8, 8, 1, 1, 11, 2, 0) op_769 (v125[7:0], v74[7:0], v769[10:0]); // 1.0
    wire [17:0] v770; shift_adder #(8, 9, 1, 1, 18, -9, 1) op_770 (v64[7:0], v128[8:0], v770[17:0]); // 2.0
    wire [12:0] v771; shift_adder #(11, 10, 1, 1, 13, 2, 0) op_771 (v129[10:0], v130[9:0], v771[12:0]); // 2.0
    wire [10:0] v772; shift_adder #(8, 11, 1, 1, 11, 0, 1) op_772 (v72[7:0], v132[10:0], v772[10:0]); // 2.0
    wire [16:0] v773; shift_adder #(11, 11, 1, 1, 17, -6, 1) op_773 (v134[10:0], v135[10:0], v773[16:0]); // 2.0
    wire [21:0] v774; shift_adder #(11, 12, 1, 1, 22, 10, 1) op_774 (v136[10:0], v137[11:0], v774[21:0]); // 2.0
    wire [11:0] v775; shift_adder #(9, 11, 1, 1, 12, -1, 0) op_775 (v138[8:0], v139[10:0], v775[11:0]); // 2.0
    wire [18:0] v776; shift_adder #(11, 11, 1, 1, 19, 8, 1) op_776 (v141[10:0], v135[10:0], v776[18:0]); // 2.0
    wire [20:0] v777; shift_adder #(11, 17, 1, 1, 21, -10, 1) op_777 (v142[10:0], v143[16:0], v777[20:0]); // 2.0
    wire [15:0] v778; shift_adder #(11, 11, 1, 1, 16, 5, 1) op_778 (v144[10:0], v145[10:0], v778[15:0]); // 2.0
    wire [14:0] v779; shift_adder #(11, 11, 1, 1, 15, -4, 1) op_779 (v147[10:0], v148[10:0], v779[14:0]); // 2.0
    wire [23:0] v780; shift_adder #(11, 12, 1, 1, 24, 12, 1) op_780 (v150[10:0], v151[11:0], v780[23:0]); // 2.0
    wire [14:0] v781; shift_adder #(11, 11, 1, 1, 15, 4, 0) op_781 (v153[10:0], v154[10:0], v781[14:0]); // 2.0
    wire [18:0] v782; shift_adder #(11, 11, 1, 1, 19, -8, 1) op_782 (v155[10:0], v156[10:0], v782[18:0]); // 2.0
    wire [16:0] v783; shift_adder #(11, 11, 1, 1, 17, -6, 1) op_783 (v157[10:0], v158[10:0], v783[16:0]); // 2.0
    wire [24:0] v784; shift_adder #(12, 25, 1, 1, 25, -9, 0) op_784 (v159[11:0], v160[24:0], v784[24:0]); // 2.0
    wire [10:0] v785; shift_adder #(8, 11, 1, 1, 11, -1, 1) op_785 (v90[7:0], v162[10:0], v785[10:0]); // 2.0
    wire [13:0] v786; shift_adder #(11, 12, 1, 1, 14, -3, 0) op_786 (v163[10:0], v164[11:0], v786[13:0]); // 2.0
    wire [13:0] v787; shift_adder #(8, 11, 1, 1, 14, -5, 1) op_787 (v78[7:0], v165[10:0], v787[13:0]); // 2.0
    wire [22:0] v788; shift_adder #(16, 18, 1, 1, 23, 5, 1) op_788 (v166[15:0], v167[17:0], v788[22:0]); // 2.0
    wire [17:0] v789; shift_adder #(11, 11, 1, 1, 18, -7, 0) op_789 (v168[10:0], v169[10:0], v789[17:0]); // 2.0
    wire [12:0] v790; shift_adder #(8, 11, 1, 1, 13, 2, 1) op_790 (v107[7:0], v171[10:0], v790[12:0]); // 2.0
    wire [24:0] v791; shift_adder #(8, 11, 1, 1, 25, 14, 1) op_791 (v92[7:0], v172[10:0], v791[24:0]); // 2.0
    wire [12:0] v792; shift_adder #(8, 11, 1, 1, 13, 2, 1) op_792 (v75[7:0], v173[10:0], v792[12:0]); // 2.0
    wire [12:0] v793; shift_adder #(8, 11, 1, 1, 13, 2, 1) op_793 (v110[7:0], v175[10:0], v793[12:0]); // 2.0
    wire [11:0] v794; shift_adder #(8, 11, 1, 1, 12, -2, 1) op_794 (v80[7:0], v177[10:0], v794[11:0]); // 2.0
    wire [12:0] v795; shift_adder #(11, 11, 1, 1, 13, 2, 1) op_795 (v141[10:0], v178[10:0], v795[12:0]); // 2.0
    wire [24:0] v796; shift_adder #(11, 12, 1, 1, 25, -14, 0) op_796 (v179[10:0], v180[11:0], v796[24:0]); // 2.0
    wire [11:0] v797; shift_adder #(11, 11, 1, 1, 12, -1, 1) op_797 (v181[10:0], v182[10:0], v797[11:0]); // 2.0
    wire [26:0] v798; shift_adder #(12, 12, 1, 1, 27, 15, 0) op_798 (v183[11:0], v184[11:0], v798[26:0]); // 2.0
    wire [13:0] v799; shift_adder #(8, 11, 1, 1, 14, 3, 0) op_799 (v114[7:0], v185[10:0], v799[13:0]); // 2.0
    wire [12:0] v800; shift_adder #(12, 11, 1, 1, 13, 1, 0) op_800 (v186[11:0], v187[10:0], v800[12:0]); // 2.0
    wire [11:0] v801; shift_adder #(11, 11, 1, 1, 12, 1, 1) op_801 (v188[10:0], v141[10:0], v801[11:0]); // 2.0
    wire [25:0] v802; shift_adder #(8, 11, 1, 1, 26, -17, 0) op_802 (v83[7:0], v190[10:0], v802[25:0]); // 2.0
    wire [12:0] v803; shift_adder #(8, 11, 1, 1, 13, -4, 0) op_803 (v118[7:0], v193[10:0], v803[12:0]); // 2.0
    wire [21:0] v804; shift_adder #(8, 12, 1, 1, 22, 10, 0) op_804 (v109[7:0], v194[11:0], v804[21:0]); // 2.0
    wire [18:0] v805; shift_adder #(11, 11, 1, 1, 19, -8, 0) op_805 (v148[10:0], v195[10:0], v805[18:0]); // 2.0
    wire [19:0] v806; shift_adder #(19, 11, 1, 1, 20, 8, 0) op_806 (v196[18:0], v152[10:0], v806[19:0]); // 2.0
    wire [13:0] v807; shift_adder #(11, 13, 1, 1, 14, 1, 1) op_807 (v197[10:0], v198[12:0], v807[13:0]); // 2.0
    wire [11:0] v808; shift_adder #(11, 11, 1, 1, 12, -1, 1) op_808 (v200[10:0], v201[10:0], v808[11:0]); // 2.0
    wire [19:0] v809; shift_adder #(11, 12, 1, 1, 20, -9, 0) op_809 (v131[10:0], v202[11:0], v809[19:0]); // 2.0
    wire [25:0] v810; shift_adder #(11, 12, 1, 1, 26, -15, 1) op_810 (v203[10:0], v204[11:0], v810[25:0]); // 2.0
    wire [22:0] v811; shift_adder #(8, 12, 1, 1, 23, 11, 0) op_811 (v94[7:0], v205[11:0], v811[22:0]); // 2.0
    wire [28:0] v812; shift_adder #(8, 11, 1, 1, 29, 18, 1) op_812 (v84[7:0], v203[10:0], v812[28:0]); // 2.0
    wire [12:0] v813; shift_adder #(8, 11, 1, 1, 13, 2, 1) op_813 (v99[7:0], v206[10:0], v813[12:0]); // 2.0
    wire [15:0] v814; shift_adder #(11, 12, 1, 1, 16, 4, 1) op_814 (v150[10:0], v207[11:0], v814[15:0]); // 2.0
    wire [14:0] v815; shift_adder #(11, 11, 1, 1, 15, 4, 0) op_815 (v199[10:0], v208[10:0], v815[14:0]); // 2.0
    wire [17:0] v816; shift_adder #(11, 11, 1, 1, 18, -7, 0) op_816 (v209[10:0], v210[10:0], v816[17:0]); // 2.0
    wire [12:0] v817; shift_adder #(11, 11, 1, 1, 13, 2, 1) op_817 (v211[10:0], v212[10:0], v817[12:0]); // 2.0
    wire [12:0] v818; shift_adder #(11, 12, 1, 1, 13, -2, 0) op_818 (v213[10:0], v214[11:0], v818[12:0]); // 2.0
    wire [16:0] v819; shift_adder #(11, 11, 1, 1, 17, -6, 0) op_819 (v216[10:0], v217[10:0], v819[16:0]); // 2.0
    wire [11:0] v820; shift_adder #(11, 11, 1, 1, 12, 0, 1) op_820 (v218[10:0], v219[10:0], v820[11:0]); // 2.0
    wire [10:0] v821; shift_adder #(8, 11, 1, 1, 11, -1, 0) op_821 (v71[7:0], v203[10:0], v821[10:0]); // 2.0
    wire [10:0] v822; shift_adder #(9, 10, 1, 1, 11, 0, 0) op_822 (v221[8:0], v222[9:0], v822[10:0]); // 2.0
    wire [12:0] v823; shift_adder #(11, 12, 1, 1, 13, -1, 0) op_823 (v223[10:0], v224[11:0], v823[12:0]); // 2.0
    wire [11:0] v824; shift_adder #(11, 11, 1, 1, 12, 1, 1) op_824 (v152[10:0], v185[10:0], v824[11:0]); // 2.0
    wire [11:0] v825; shift_adder #(8, 11, 1, 1, 12, 1, 0) op_825 (v69[7:0], v171[10:0], v825[11:0]); // 2.0
    wire [12:0] v826; shift_adder #(8, 11, 1, 1, 13, 2, 1) op_826 (v94[7:0], v208[10:0], v826[12:0]); // 2.0
    wire [13:0] v827; shift_adder #(10, 14, 1, 1, 14, 0, 0) op_827 (v225[9:0], v226[13:0], v827[13:0]); // 2.0
    wire [12:0] v828; shift_adder #(8, 11, 1, 1, 13, -4, 1) op_828 (v77[7:0], v161[10:0], v828[12:0]); // 2.0
    wire [24:0] v829; shift_adder #(8, 12, 1, 1, 25, -16, 0) op_829 (v111[7:0], v227[11:0], v829[24:0]); // 2.0
    wire [13:0] v830; shift_adder #(8, 11, 1, 1, 14, -5, 1) op_830 (v69[7:0], v229[10:0], v830[13:0]); // 2.0
    wire [11:0] v831; shift_adder #(9, 9, 1, 1, 12, -2, 0) op_831 (v230[8:0], v231[8:0], v831[11:0]); // 2.0
    wire [16:0] v832; shift_adder #(11, 12, 1, 1, 17, 5, 1) op_832 (v233[10:0], v224[11:0], v832[16:0]); // 2.0
    wire [12:0] v833; shift_adder #(8, 11, 1, 1, 13, 2, 1) op_833 (v101[7:0], v234[10:0], v833[12:0]); // 2.0
    wire [12:0] v834; shift_adder #(11, 11, 1, 1, 13, -2, 0) op_834 (v237[10:0], v238[10:0], v834[12:0]); // 2.0
    wire [11:0] v835; shift_adder #(8, 11, 1, 1, 12, -3, 1) op_835 (v122[7:0], v237[10:0], v835[11:0]); // 2.0
    wire [15:0] v836; shift_adder #(12, 16, 1, 1, 16, -2, 0) op_836 (v239[11:0], v240[15:0], v836[15:0]); // 2.0
    wire [12:0] v837; shift_adder #(8, 11, 1, 1, 13, -4, 0) op_837 (v127[7:0], v241[10:0], v837[12:0]); // 2.0
    wire [26:0] v838; shift_adder #(11, 11, 1, 1, 27, -16, 0) op_838 (v139[10:0], v242[10:0], v838[26:0]); // 2.0
    wire [14:0] v839; shift_adder #(11, 11, 1, 1, 15, -4, 0) op_839 (v244[10:0], v244[10:0], v839[14:0]); // 2.0
    wire [14:0] v840; shift_adder #(11, 11, 1, 1, 15, 4, 0) op_840 (v245[10:0], v233[10:0], v840[14:0]); // 2.0
    wire [19:0] v841; shift_adder #(11, 11, 1, 1, 20, -9, 0) op_841 (v133[10:0], v246[10:0], v841[19:0]); // 2.0
    wire [13:0] v842; shift_adder #(8, 11, 1, 1, 14, -5, 1) op_842 (v84[7:0], v200[10:0], v842[13:0]); // 2.0
    wire [11:0] v843; shift_adder #(11, 10, 1, 1, 12, 1, 0) op_843 (v187[10:0], v248[9:0], v843[11:0]); // 2.0
    wire [21:0] v844; shift_adder #(11, 14, 1, 1, 22, -11, 1) op_844 (v199[10:0], v249[13:0], v844[21:0]); // 2.0
    wire [12:0] v845; shift_adder #(8, 11, 1, 1, 13, 2, 1) op_845 (v119[7:0], v250[10:0], v845[12:0]); // 2.0
    wire [10:0] v846; shift_adder #(8, 11, 1, 1, 11, -1, 0) op_846 (v111[7:0], v251[10:0], v846[10:0]); // 2.0
    wire [16:0] v847; shift_adder #(15, 10, 1, 1, 17, 7, 0) op_847 (v253[14:0], v254[9:0], v847[16:0]); // 2.0
    wire [11:0] v848; shift_adder #(8, 11, 1, 1, 12, -2, 0) op_848 (v82[7:0], v203[10:0], v848[11:0]); // 2.0
    wire [15:0] v849; shift_adder #(11, 11, 1, 1, 16, -5, 0) op_849 (v157[10:0], v255[10:0], v849[15:0]); // 2.0
    wire [28:0] v850; shift_adder #(8, 9, 1, 1, 29, 20, 1) op_850 (v86[7:0], v256[8:0], v850[28:0]); // 2.0
    wire [22:0] v851; shift_adder #(12, 23, 1, 1, 23, -9, 0) op_851 (v257[11:0], v258[22:0], v851[22:0]); // 2.0
    wire [16:0] v852; shift_adder #(8, 11, 1, 1, 17, -8, 1) op_852 (v124[7:0], v131[10:0], v852[16:0]); // 2.0
    wire [17:0] v853; shift_adder #(11, 11, 1, 1, 18, 7, 1) op_853 (v237[10:0], v259[10:0], v853[17:0]); // 2.0
    wire [11:0] v854; shift_adder #(8, 11, 1, 1, 12, -3, 0) op_854 (v76[7:0], v171[10:0], v854[11:0]); // 2.0
    wire [10:0] v855; shift_adder #(8, 9, 1, 1, 11, -2, 1) op_855 (v79[7:0], v221[8:0], v855[10:0]); // 2.0
    wire [17:0] v856; shift_adder #(17, 10, 1, 1, 18, 7, 0) op_856 (v143[16:0], v260[9:0], v856[17:0]); // 2.0
    wire [11:0] v857; shift_adder #(11, 11, 1, 1, 12, 0, 0) op_857 (v132[10:0], v172[10:0], v857[11:0]); // 2.0
    wire [32:0] v858; shift_adder #(25, 32, 1, 1, 33, -8, 0) op_858 (v261[24:0], v262[31:0], v858[32:0]); // 2.0
    wire [12:0] v859; shift_adder #(8, 11, 1, 1, 13, 2, 1) op_859 (v114[7:0], v228[10:0], v859[12:0]); // 2.0
    wire [12:0] v860; shift_adder #(11, 12, 1, 1, 13, -1, 1) op_860 (v264[10:0], v265[11:0], v860[12:0]); // 2.0
    wire [12:0] v861; shift_adder #(11, 12, 1, 1, 13, -1, 0) op_861 (v266[10:0], v267[11:0], v861[12:0]); // 2.0
    wire [11:0] v862; shift_adder #(11, 11, 1, 1, 12, 0, 1) op_862 (v190[10:0], v150[10:0], v862[11:0]); // 2.0
    wire [11:0] v863; shift_adder #(8, 11, 1, 1, 12, -3, 0) op_863 (v99[7:0], v223[10:0], v863[11:0]); // 2.0
    wire [23:0] v864; shift_adder #(11, 11, 1, 1, 24, 13, 0) op_864 (v238[10:0], v195[10:0], v864[23:0]); // 2.0
    wire [17:0] v865; shift_adder #(8, 11, 1, 1, 18, 7, 0) op_865 (v107[7:0], v269[10:0], v865[17:0]); // 2.0
    wire [14:0] v866; shift_adder #(8, 11, 1, 1, 15, 4, 1) op_866 (v77[7:0], v244[10:0], v866[14:0]); // 2.0
    wire [11:0] v867; shift_adder #(11, 11, 1, 1, 12, 0, 0) op_867 (v175[10:0], v270[10:0], v867[11:0]); // 2.0
    wire [21:0] v868; shift_adder #(13, 10, 1, 1, 22, -9, 0) op_868 (v272[12:0], v273[9:0], v868[21:0]); // 2.0
    wire [16:0] v869; shift_adder #(11, 12, 1, 1, 17, -6, 0) op_869 (v274[10:0], v224[11:0], v869[16:0]); // 2.0
    wire [10:0] v870; shift_adder #(8, 11, 1, 1, 11, 0, 1) op_870 (v69[7:0], v172[10:0], v870[10:0]); // 2.0
    wire [13:0] v871; shift_adder #(11, 11, 1, 1, 14, 3, 1) op_871 (v219[10:0], v275[10:0], v871[13:0]); // 2.0
    wire [17:0] v872; shift_adder #(11, 11, 1, 1, 18, 7, 0) op_872 (v144[10:0], v264[10:0], v872[17:0]); // 2.0
    wire [11:0] v873; shift_adder #(8, 11, 1, 1, 12, -3, 1) op_873 (v100[7:0], v187[10:0], v873[11:0]); // 2.0
    wire [17:0] v874; shift_adder #(11, 11, 1, 1, 18, -7, 0) op_874 (v276[10:0], v277[10:0], v874[17:0]); // 2.0
    wire [16:0] v875; shift_adder #(13, 12, 1, 1, 17, -4, 0) op_875 (v278[12:0], v279[11:0], v875[16:0]); // 2.0
    wire [16:0] v876; shift_adder #(11, 11, 1, 1, 17, 6, 0) op_876 (v206[10:0], v211[10:0], v876[16:0]); // 2.0
    wire [12:0] v877; shift_adder #(12, 11, 1, 1, 13, 2, 1) op_877 (v280[11:0], v281[10:0], v877[12:0]); // 2.0
    wire [13:0] v878; shift_adder #(11, 10, 1, 1, 14, 4, 0) op_878 (v139[10:0], v282[9:0], v878[13:0]); // 2.0
    wire [11:0] v879; shift_adder #(11, 11, 1, 1, 12, 0, 1) op_879 (v283[10:0], v284[10:0], v879[11:0]); // 2.0
    wire [12:0] v880; shift_adder #(8, 11, 1, 1, 13, 2, 1) op_880 (v124[7:0], v218[10:0], v880[12:0]); // 2.0
    wire [16:0] v881; shift_adder #(11, 11, 1, 1, 17, -6, 1) op_881 (v140[10:0], v287[10:0], v881[16:0]); // 2.0
    wire [12:0] v882; shift_adder #(8, 11, 1, 1, 13, -4, 0) op_882 (v95[7:0], v289[10:0], v882[12:0]); // 2.0
    wire [12:0] v883; shift_adder #(8, 11, 1, 1, 13, -4, 1) op_883 (v127[7:0], v241[10:0], v883[12:0]); // 2.0
    wire [12:0] v884; shift_adder #(8, 11, 1, 1, 13, 2, 1) op_884 (v125[7:0], v276[10:0], v884[12:0]); // 2.0
    wire [10:0] v885; shift_adder #(8, 11, 1, 1, 11, -1, 0) op_885 (v89[7:0], v244[10:0], v885[10:0]); // 2.0
    wire [14:0] v886; shift_adder #(12, 11, 1, 1, 15, -3, 0) op_886 (v292[11:0], v293[10:0], v886[14:0]); // 2.0
    wire [16:0] v887; shift_adder #(11, 11, 1, 1, 17, 6, 1) op_887 (v210[10:0], v294[10:0], v887[16:0]); // 2.0
    wire [12:0] v888; shift_adder #(13, 11, 1, 1, 13, 1, 0) op_888 (v296[12:0], v255[10:0], v888[12:0]); // 2.0
    wire [16:0] v889; shift_adder #(11, 12, 1, 1, 17, 5, 1) op_889 (v218[10:0], v243[11:0], v889[16:0]); // 2.0
    wire [16:0] v890; shift_adder #(11, 11, 1, 1, 17, 6, 0) op_890 (v156[10:0], v297[10:0], v890[16:0]); // 2.0
    wire [12:0] v891; shift_adder #(11, 11, 1, 1, 13, -2, 1) op_891 (v218[10:0], v136[10:0], v891[12:0]); // 2.0
    wire [12:0] v892; shift_adder #(11, 11, 1, 1, 13, -2, 1) op_892 (v283[10:0], v211[10:0], v892[12:0]); // 2.0
    wire [14:0] v893; shift_adder #(8, 11, 1, 1, 15, 4, 0) op_893 (v95[7:0], v193[10:0], v893[14:0]); // 2.0
    wire [14:0] v894; shift_adder #(12, 12, 1, 1, 15, 3, 0) op_894 (v183[11:0], v204[11:0], v894[14:0]); // 2.0
    wire [16:0] v895; shift_adder #(11, 11, 1, 1, 17, -6, 0) op_895 (v298[10:0], v299[10:0], v895[16:0]); // 2.0
    wire [11:0] v896; shift_adder #(11, 11, 1, 1, 12, -1, 0) op_896 (v140[10:0], v299[10:0], v896[11:0]); // 2.0
    wire [16:0] v897; shift_adder #(11, 11, 1, 1, 17, -6, 0) op_897 (v199[10:0], v161[10:0], v897[16:0]); // 2.0
    wire [12:0] v898; shift_adder #(11, 11, 1, 1, 13, -2, 1) op_898 (v300[10:0], v213[10:0], v898[12:0]); // 2.0
    wire [13:0] v899; shift_adder #(11, 11, 1, 1, 14, 3, 1) op_899 (v145[10:0], v150[10:0], v899[13:0]); // 2.0
    wire [12:0] v900; shift_adder #(11, 11, 1, 1, 13, -2, 1) op_900 (v219[10:0], v195[10:0], v900[12:0]); // 2.0
    wire [15:0] v901; shift_adder #(8, 11, 1, 1, 16, 5, 0) op_901 (v67[7:0], v283[10:0], v901[15:0]); // 2.0
    wire [14:0] v902; shift_adder #(11, 11, 1, 1, 15, 4, 1) op_902 (v242[10:0], v287[10:0], v902[14:0]); // 2.0
    wire [18:0] v903; shift_adder #(11, 9, 1, 1, 19, 9, 0) op_903 (v301[10:0], v302[8:0], v903[18:0]); // 2.0
    wire [14:0] v904; shift_adder #(11, 11, 1, 1, 15, 4, 0) op_904 (v215[10:0], v266[10:0], v904[14:0]); // 2.0
    wire [14:0] v905; shift_adder #(11, 11, 1, 1, 15, 4, 1) op_905 (v201[10:0], v303[10:0], v905[14:0]); // 2.0
    wire [21:0] v906; shift_adder #(8, 11, 1, 1, 22, 11, 0) op_906 (v68[7:0], v223[10:0], v906[21:0]); // 2.0
    wire [20:0] v907; shift_adder #(8, 11, 1, 1, 21, 10, 0) op_907 (v88[7:0], v209[10:0], v907[20:0]); // 2.0
    wire [21:0] v908; shift_adder #(12, 12, 1, 1, 22, 10, 1) op_908 (v304[11:0], v305[11:0], v908[21:0]); // 2.0
    wire [21:0] v909; shift_adder #(8, 11, 1, 1, 22, 11, 1) op_909 (v84[7:0], v188[10:0], v909[21:0]); // 2.0
    wire [18:0] v910; shift_adder #(17, 10, 1, 1, 19, 9, 0) op_910 (v306[16:0], v307[9:0], v910[18:0]); // 2.0
    wire [18:0] v911; shift_adder #(12, 15, 1, 1, 19, -7, 1) op_911 (v285[11:0], v308[14:0], v911[18:0]); // 2.0
    wire [26:0] v912; shift_adder #(9, 20, 1, 1, 27, -17, 1) op_912 (v309[8:0], v310[19:0], v912[26:0]); // 2.0
    wire [14:0] v913; shift_adder #(11, 11, 1, 1, 15, -4, 1) op_913 (v141[10:0], v135[10:0], v913[14:0]); // 2.0
    wire [14:0] v914; shift_adder #(8, 10, 1, 1, 15, -6, 1) op_914 (v91[7:0], v311[9:0], v914[14:0]); // 2.0
    wire [12:0] v915; shift_adder #(8, 11, 1, 1, 13, 2, 1) op_915 (v82[7:0], v140[10:0], v915[12:0]); // 2.0
    wire [24:0] v916; shift_adder #(8, 11, 1, 1, 25, -16, 0) op_916 (v91[7:0], v238[10:0], v916[24:0]); // 2.0
    wire [16:0] v917; shift_adder #(11, 12, 1, 1, 17, 5, 1) op_917 (v213[10:0], v314[11:0], v917[16:0]); // 2.0
    wire [21:0] v918; shift_adder #(19, 9, 1, 1, 22, 12, 1) op_918 (v315[18:0], v316[8:0], v918[21:0]); // 2.0
    wire [11:0] v919; shift_adder #(11, 11, 1, 1, 12, -1, 1) op_919 (v317[10:0], v200[10:0], v919[11:0]); // 2.0
    wire [12:0] v920; shift_adder #(8, 11, 1, 1, 13, 2, 1) op_920 (v71[7:0], v131[10:0], v920[12:0]); // 2.0
    wire [16:0] v921; shift_adder #(8, 11, 1, 1, 17, 6, 0) op_921 (v78[7:0], v250[10:0], v921[16:0]); // 2.0
    wire [14:0] v922; shift_adder #(8, 11, 1, 1, 15, -6, 0) op_922 (v69[7:0], v269[10:0], v922[14:0]); // 2.0
    wire [12:0] v923; shift_adder #(11, 11, 1, 1, 13, 2, 1) op_923 (v275[10:0], v185[10:0], v923[12:0]); // 2.0
    wire [11:0] v924; shift_adder #(11, 11, 1, 1, 12, -1, 1) op_924 (v270[10:0], v181[10:0], v924[11:0]); // 2.0
    wire [19:0] v925; shift_adder #(11, 11, 1, 1, 20, 9, 1) op_925 (v178[10:0], v320[10:0], v925[19:0]); // 2.0
    wire [17:0] v926; shift_adder #(8, 11, 1, 1, 18, -9, 1) op_926 (v100[7:0], v233[10:0], v926[17:0]); // 2.0
    wire [15:0] v927; shift_adder #(11, 11, 1, 1, 16, -5, 1) op_927 (v148[10:0], v148[10:0], v927[15:0]); // 2.0
    wire [13:0] v928; shift_adder #(11, 12, 1, 1, 14, -3, 0) op_928 (v195[10:0], v321[11:0], v928[13:0]); // 2.0
    wire [11:0] v929; shift_adder #(8, 9, 1, 1, 12, 2, 1) op_929 (v123[7:0], v322[8:0], v929[11:0]); // 2.0
    wire [26:0] v930; shift_adder #(11, 11, 1, 1, 27, 16, 1) op_930 (v323[10:0], v161[10:0], v930[26:0]); // 2.0
    wire [18:0] v931; shift_adder #(12, 11, 1, 1, 19, -7, 1) op_931 (v174[11:0], v191[10:0], v931[18:0]); // 2.0
    wire [12:0] v932; shift_adder #(8, 11, 1, 1, 13, 2, 1) op_932 (v106[7:0], v223[10:0], v932[12:0]); // 2.0
    wire [26:0] v933; shift_adder #(11, 11, 1, 1, 27, -16, 1) op_933 (v251[10:0], v200[10:0], v933[26:0]); // 2.0
    wire [11:0] v934; shift_adder #(11, 11, 1, 1, 12, 1, 0) op_934 (v132[10:0], v324[10:0], v934[11:0]); // 2.0
    wire [11:0] v935; shift_adder #(11, 11, 1, 1, 12, 1, 0) op_935 (v237[10:0], v275[10:0], v935[11:0]); // 2.0
    wire [11:0] v936; shift_adder #(11, 11, 1, 1, 12, 0, 1) op_936 (v238[10:0], v223[10:0], v936[11:0]); // 2.0
    wire [13:0] v937; shift_adder #(12, 13, 1, 1, 14, 1, 0) op_937 (v325[11:0], v326[12:0], v937[13:0]); // 2.0
    wire [17:0] v938; shift_adder #(11, 11, 1, 1, 18, 7, 1) op_938 (v244[10:0], v294[10:0], v938[17:0]); // 2.0
    wire [17:0] v939; shift_adder #(8, 13, 1, 1, 18, -9, 0) op_939 (v121[7:0], v327[12:0], v939[17:0]); // 2.0
    wire [17:0] v940; shift_adder #(8, 11, 1, 1, 18, -9, 0) op_940 (v82[7:0], v328[10:0], v940[17:0]); // 2.0
    wire [10:0] v941; shift_adder #(8, 11, 1, 1, 11, 0, 1) op_941 (v67[7:0], v329[10:0], v941[10:0]); // 2.0
    wire [11:0] v942; shift_adder #(11, 11, 1, 1, 12, 0, 0) op_942 (v152[10:0], v300[10:0], v942[11:0]); // 2.0
    wire [20:0] v943; shift_adder #(11, 11, 1, 1, 21, -10, 0) op_943 (v144[10:0], v193[10:0], v943[20:0]); // 2.0
    wire [18:0] v944; shift_adder #(8, 11, 1, 1, 19, -10, 1) op_944 (v86[7:0], v147[10:0], v944[18:0]); // 2.0
    wire [14:0] v945; shift_adder #(11, 11, 1, 1, 15, -4, 1) op_945 (v178[10:0], v319[10:0], v945[14:0]); // 2.0
    wire [15:0] v946; shift_adder #(8, 11, 1, 1, 16, 5, 0) op_946 (v97[7:0], v210[10:0], v946[15:0]); // 2.0
    wire [31:0] v947; shift_adder #(10, 32, 1, 1, 32, -21, 0) op_947 (v331[9:0], v332[31:0], v947[31:0]); // 2.0
    wire [12:0] v948; shift_adder #(11, 11, 1, 1, 13, 2, 0) op_948 (v153[10:0], v334[10:0], v948[12:0]); // 2.0
    wire [17:0] v949; shift_adder #(11, 17, 1, 1, 18, 1, 1) op_949 (v199[10:0], v335[16:0], v949[17:0]); // 2.0
    wire [13:0] v950; shift_adder #(12, 12, 1, 1, 14, 2, 1) op_950 (v336[11:0], v337[11:0], v950[13:0]); // 2.0
    wire [20:0] v951; shift_adder #(11, 11, 1, 1, 21, 10, 1) op_951 (v210[10:0], v139[10:0], v951[20:0]); // 2.0
    wire [16:0] v952; shift_adder #(11, 11, 1, 1, 17, -6, 0) op_952 (v171[10:0], v338[10:0], v952[16:0]); // 2.0
    wire [12:0] v953; shift_adder #(12, 11, 1, 1, 13, 1, 0) op_953 (v339[11:0], v148[10:0], v953[12:0]); // 2.0
    wire [10:0] v954; shift_adder #(8, 11, 1, 1, 11, 0, 1) op_954 (v113[7:0], v158[10:0], v954[10:0]); // 2.0
    wire [33:0] v955; shift_adder #(9, 10, 1, 1, 34, -24, 1) op_955 (v340[8:0], v307[9:0], v955[33:0]); // 2.0
    wire [11:0] v956; shift_adder #(11, 11, 1, 1, 12, -1, 0) op_956 (v264[10:0], v341[10:0], v956[11:0]); // 2.0
    wire [11:0] v957; shift_adder #(11, 11, 1, 1, 12, 0, 0) op_957 (v176[10:0], v188[10:0], v957[11:0]); // 2.0
    wire [13:0] v958; shift_adder #(11, 14, 1, 1, 14, -2, 0) op_958 (v269[10:0], v342[13:0], v958[13:0]); // 2.0
    wire [15:0] v959; shift_adder #(11, 11, 1, 1, 16, -5, 1) op_959 (v250[10:0], v276[10:0], v959[15:0]); // 2.0
    wire [13:0] v960; shift_adder #(11, 13, 1, 1, 14, -3, 0) op_960 (v343[10:0], v344[12:0], v960[13:0]); // 2.0
    wire [10:0] v961; shift_adder #(8, 11, 1, 1, 11, 0, 0) op_961 (v94[7:0], v345[10:0], v961[10:0]); // 2.0
    wire [10:0] v962; shift_adder #(8, 11, 1, 1, 11, 0, 0) op_962 (v77[7:0], v173[10:0], v962[10:0]); // 2.0
    wire [16:0] v963; shift_adder #(8, 12, 1, 1, 17, 5, 1) op_963 (v119[7:0], v347[11:0], v963[16:0]); // 2.0
    wire [13:0] v964; shift_adder #(8, 11, 1, 1, 14, -5, 0) op_964 (v100[7:0], v217[10:0], v964[13:0]); // 2.0
    wire [11:0] v965; shift_adder #(8, 9, 1, 1, 12, -3, 0) op_965 (v123[7:0], v302[8:0], v965[11:0]); // 2.0
    wire [16:0] v966; shift_adder #(17, 13, 1, 1, 17, 1, 0) op_966 (v348[16:0], v349[12:0], v966[16:0]); // 2.0
    wire [16:0] v967; shift_adder #(8, 16, 1, 1, 17, 1, 1) op_967 (v99[7:0], v350[15:0], v967[16:0]); // 2.0
    wire [17:0] v968; shift_adder #(11, 11, 1, 1, 18, 7, 1) op_968 (v203[10:0], v157[10:0], v968[17:0]); // 2.0
    wire [14:0] v969; shift_adder #(11, 11, 1, 1, 15, -4, 1) op_969 (v163[10:0], v352[10:0], v969[14:0]); // 2.0
    wire [15:0] v970; shift_adder #(8, 11, 1, 1, 16, 5, 1) op_970 (v118[7:0], v241[10:0], v970[15:0]); // 2.0
    wire [11:0] v971; shift_adder #(11, 11, 1, 1, 12, 0, 1) op_971 (v208[10:0], v352[10:0], v971[11:0]); // 2.0
    wire [16:0] v972; shift_adder #(11, 11, 1, 1, 17, 6, 0) op_972 (v215[10:0], v338[10:0], v972[16:0]); // 2.0
    wire [11:0] v973; shift_adder #(11, 11, 1, 1, 12, 0, 1) op_973 (v134[10:0], v353[10:0], v973[11:0]); // 2.0
    wire [12:0] v974; shift_adder #(11, 12, 1, 1, 13, 1, 0) op_974 (v297[10:0], v354[11:0], v974[12:0]); // 2.0
    wire [13:0] v975; shift_adder #(8, 11, 1, 1, 14, 3, 0) op_975 (v86[7:0], v270[10:0], v975[13:0]); // 2.0
    wire [13:0] v976; shift_adder #(11, 11, 1, 1, 14, 3, 0) op_976 (v175[10:0], v320[10:0], v976[13:0]); // 2.0
    wire [17:0] v977; shift_adder #(11, 18, 1, 1, 18, -6, 1) op_977 (v276[10:0], v167[17:0], v977[17:0]); // 2.0
    wire [12:0] v978; shift_adder #(11, 12, 1, 1, 13, -2, 0) op_978 (v287[10:0], v355[11:0], v978[12:0]); // 2.0
    wire [25:0] v979; shift_adder #(11, 10, 1, 1, 26, -15, 0) op_979 (v298[10:0], v130[9:0], v979[25:0]); // 2.0
    wire [22:0] v980; shift_adder #(11, 23, 1, 1, 23, -11, 0) op_980 (v237[10:0], v258[22:0], v980[22:0]); // 2.0
    wire [11:0] v981; shift_adder #(11, 11, 1, 1, 12, 0, 0) op_981 (v301[10:0], v303[10:0], v981[11:0]); // 2.0
    wire [16:0] v982; shift_adder #(8, 11, 1, 1, 17, -8, 0) op_982 (v89[7:0], v152[10:0], v982[16:0]); // 2.0
    wire [12:0] v983; shift_adder #(11, 11, 1, 1, 13, 2, 0) op_983 (v182[10:0], v154[10:0], v983[12:0]); // 2.0
    wire [29:0] v984; shift_adder #(8, 9, 1, 1, 30, 21, 1) op_984 (v71[7:0], v351[8:0], v984[29:0]); // 2.0
    wire [12:0] v985; shift_adder #(8, 12, 1, 1, 13, -4, 1) op_985 (v101[7:0], v174[11:0], v985[12:0]); // 2.0
    wire [13:0] v986; shift_adder #(12, 11, 1, 1, 14, 3, 0) op_986 (v357[11:0], v358[10:0], v986[13:0]); // 2.0
    wire [10:0] v987; shift_adder #(10, 10, 1, 1, 11, 0, 0) op_987 (v130[9:0], v248[9:0], v987[10:0]); // 2.0
    wire [25:0] v988; shift_adder #(8, 13, 1, 1, 26, 13, 0) op_988 (v72[7:0], v359[12:0], v988[25:0]); // 2.0
    wire [17:0] v989; shift_adder #(11, 11, 1, 1, 18, -7, 0) op_989 (v157[10:0], v191[10:0], v989[17:0]); // 2.0
    wire [11:0] v990; shift_adder #(11, 11, 1, 1, 12, 0, 1) op_990 (v203[10:0], v334[10:0], v990[11:0]); // 2.0
    wire [11:0] v991; shift_adder #(11, 10, 1, 1, 12, -1, 0) op_991 (v238[10:0], v235[9:0], v991[11:0]); // 2.0
    wire [13:0] v992; shift_adder #(11, 11, 1, 1, 14, -3, 0) op_992 (v173[10:0], v300[10:0], v992[13:0]); // 2.0
    wire [14:0] v993; shift_adder #(11, 11, 1, 1, 15, 4, 1) op_993 (v147[10:0], v206[10:0], v993[14:0]); // 2.0
    wire [20:0] v994; shift_adder #(8, 11, 1, 1, 21, 10, 1) op_994 (v78[7:0], v284[10:0], v994[20:0]); // 2.0
    wire [12:0] v995; shift_adder #(11, 11, 1, 1, 13, 2, 1) op_995 (v141[10:0], v216[10:0], v995[12:0]); // 2.0
    wire [12:0] v996; shift_adder #(8, 11, 1, 1, 13, 2, 0) op_996 (v76[7:0], v165[10:0], v996[12:0]); // 2.0
    wire [13:0] v997; shift_adder #(13, 11, 1, 1, 14, 3, 0) op_997 (v327[12:0], v301[10:0], v997[13:0]); // 2.0
    wire [20:0] v998; shift_adder #(11, 11, 1, 1, 21, 10, 0) op_998 (v171[10:0], v323[10:0], v998[20:0]); // 2.0
    wire [11:0] v999; shift_adder #(11, 11, 1, 1, 12, 1, 1) op_999 (v212[10:0], v361[10:0], v999[11:0]); // 2.0
    wire [11:0] v1000; shift_adder #(11, 12, 1, 1, 12, 0, 0) op_1000 (v362[10:0], v363[11:0], v1000[11:0]); // 2.0
    wire [12:0] v1001; shift_adder #(8, 11, 1, 1, 13, 2, 1) op_1001 (v83[7:0], v142[10:0], v1001[12:0]); // 2.0
    wire [13:0] v1002; shift_adder #(8, 11, 1, 1, 14, -5, 0) op_1002 (v102[7:0], v156[10:0], v1002[13:0]); // 2.0
    wire [21:0] v1003; shift_adder #(21, 12, 1, 1, 22, 10, 0) op_1003 (v364[20:0], v365[11:0], v1003[21:0]); // 2.0
    wire [11:0] v1004; shift_adder #(11, 9, 1, 1, 12, -1, 1) op_1004 (v329[10:0], v368[8:0], v1004[11:0]); // 2.0
    wire [17:0] v1005; shift_adder #(11, 11, 1, 1, 18, -7, 1) op_1005 (v244[10:0], v275[10:0], v1005[17:0]); // 2.0
    wire [14:0] v1006; shift_adder #(11, 11, 1, 1, 15, 4, 1) op_1006 (v229[10:0], v208[10:0], v1006[14:0]); // 2.0
    wire [13:0] v1007; shift_adder #(8, 11, 1, 1, 14, 3, 1) op_1007 (v110[7:0], v259[10:0], v1007[13:0]); // 2.0
    wire [21:0] v1008; shift_adder #(9, 22, 1, 1, 22, -8, 0) op_1008 (v370[8:0], v371[21:0], v1008[21:0]); // 2.0
    wire [18:0] v1009; shift_adder #(11, 11, 1, 1, 19, -8, 1) op_1009 (v181[10:0], v323[10:0], v1009[18:0]); // 2.0
    wire [14:0] v1010; shift_adder #(11, 11, 1, 1, 15, -4, 1) op_1010 (v131[10:0], v131[10:0], v1010[14:0]); // 2.0
    wire [14:0] v1011; shift_adder #(8, 11, 1, 1, 15, -6, 0) op_1011 (v74[7:0], v301[10:0], v1011[14:0]); // 2.0
    wire [14:0] v1012; shift_adder #(11, 11, 1, 1, 15, 4, 1) op_1012 (v177[10:0], v284[10:0], v1012[14:0]); // 2.0
    wire [13:0] v1013; shift_adder #(11, 11, 1, 1, 14, -3, 0) op_1013 (v215[10:0], v374[10:0], v1013[13:0]); // 2.0
    wire [13:0] v1014; shift_adder #(8, 11, 1, 1, 14, 3, 0) op_1014 (v64[7:0], v375[10:0], v1014[13:0]); // 2.0
    wire [14:0] v1015; shift_adder #(11, 11, 1, 1, 15, -4, 1) op_1015 (v144[10:0], v215[10:0], v1015[14:0]); // 2.0
    wire [16:0] v1016; shift_adder #(11, 11, 1, 1, 17, -6, 1) op_1016 (v319[10:0], v246[10:0], v1016[16:0]); // 2.0
    wire [24:0] v1017; shift_adder #(18, 11, 1, 1, 25, 14, 0) op_1017 (v378[17:0], v379[10:0], v1017[24:0]); // 2.0
    wire [12:0] v1018; shift_adder #(11, 12, 1, 1, 13, -1, 0) op_1018 (v244[10:0], v380[11:0], v1018[12:0]); // 2.0
    wire [14:0] v1019; shift_adder #(11, 11, 1, 1, 15, 4, 0) op_1019 (v229[10:0], v234[10:0], v1019[14:0]); // 2.0
    wire [15:0] v1020; shift_adder #(11, 11, 1, 1, 16, 5, 0) op_1020 (v218[10:0], v375[10:0], v1020[15:0]); // 2.0
    wire [12:0] v1021; shift_adder #(8, 11, 1, 1, 13, 2, 1) op_1021 (v76[7:0], v155[10:0], v1021[12:0]); // 2.0
    wire [27:0] v1022; shift_adder #(8, 11, 1, 1, 28, -19, 0) op_1022 (v123[7:0], v251[10:0], v1022[27:0]); // 2.0
    wire [16:0] v1023; shift_adder #(8, 11, 1, 1, 17, -8, 1) op_1023 (v115[7:0], v361[10:0], v1023[16:0]); // 2.0
    wire [12:0] v1024; shift_adder #(8, 11, 1, 1, 13, -4, 1) op_1024 (v83[7:0], v144[10:0], v1024[12:0]); // 2.0
    wire [11:0] v1025; shift_adder #(11, 11, 1, 1, 12, 1, 1) op_1025 (v238[10:0], v154[10:0], v1025[11:0]); // 2.0
    wire [12:0] v1026; shift_adder #(11, 11, 1, 1, 13, 2, 1) op_1026 (v141[10:0], v266[10:0], v1026[12:0]); // 2.0
    wire [14:0] v1027; shift_adder #(11, 11, 1, 1, 15, -4, 1) op_1027 (v182[10:0], v187[10:0], v1027[14:0]); // 2.0
    wire [15:0] v1028; shift_adder #(16, 12, 1, 1, 16, 0, 0) op_1028 (v166[15:0], v382[11:0], v1028[15:0]); // 2.0
    wire [12:0] v1029; shift_adder #(8, 11, 1, 1, 13, -4, 1) op_1029 (v88[7:0], v188[10:0], v1029[12:0]); // 2.0
    wire [12:0] v1030; shift_adder #(8, 11, 1, 1, 13, -4, 0) op_1030 (v120[7:0], v203[10:0], v1030[12:0]); // 2.0
    wire [11:0] v1031; shift_adder #(11, 11, 1, 1, 12, 0, 0) op_1031 (v177[10:0], v201[10:0], v1031[11:0]); // 2.0
    wire [17:0] v1032; shift_adder #(11, 11, 1, 1, 18, -7, 0) op_1032 (v223[10:0], v269[10:0], v1032[17:0]); // 2.0
    wire [15:0] v1033; shift_adder #(9, 12, 1, 1, 16, -6, 0) op_1033 (v384[8:0], v385[11:0], v1033[15:0]); // 2.0
    wire [12:0] v1034; shift_adder #(8, 11, 1, 1, 13, 2, 1) op_1034 (v123[7:0], v219[10:0], v1034[12:0]); // 2.0
    wire [11:0] v1035; shift_adder #(11, 11, 1, 1, 12, 1, 0) op_1035 (v216[10:0], v169[10:0], v1035[11:0]); // 2.0
    wire [18:0] v1036; shift_adder #(11, 11, 1, 1, 19, 8, 0) op_1036 (v153[10:0], v324[10:0], v1036[18:0]); // 2.0
    wire [16:0] v1037; shift_adder #(8, 12, 1, 1, 17, -8, 0) op_1037 (v90[7:0], v265[11:0], v1037[16:0]); // 2.0
    wire [14:0] v1038; shift_adder #(8, 11, 1, 1, 15, -6, 1) op_1038 (v87[7:0], v200[10:0], v1038[14:0]); // 2.0
    wire [13:0] v1039; shift_adder #(11, 11, 1, 1, 14, 3, 1) op_1039 (v237[10:0], v367[10:0], v1039[13:0]); // 2.0
    wire [20:0] v1040; shift_adder #(11, 11, 1, 1, 21, 10, 1) op_1040 (v386[10:0], v259[10:0], v1040[20:0]); // 2.0
    wire [12:0] v1041; shift_adder #(8, 11, 1, 1, 13, -4, 1) op_1041 (v67[7:0], v362[10:0], v1041[12:0]); // 2.0
    wire [25:0] v1042; shift_adder #(12, 12, 1, 1, 26, 14, 0) op_1042 (v387[11:0], v383[11:0], v1042[25:0]); // 2.0
    wire [11:0] v1043; shift_adder #(11, 11, 1, 1, 12, 0, 1) op_1043 (v175[10:0], v270[10:0], v1043[11:0]); // 2.0
    wire [23:0] v1044; shift_adder #(11, 11, 1, 1, 24, 13, 0) op_1044 (v276[10:0], v190[10:0], v1044[23:0]); // 2.0
    wire [13:0] v1045; shift_adder #(11, 12, 1, 1, 14, -3, 1) op_1045 (v299[10:0], v388[11:0], v1045[13:0]); // 2.0
    wire [12:0] v1046; shift_adder #(8, 11, 1, 1, 13, -4, 1) op_1046 (v120[7:0], v132[10:0], v1046[12:0]); // 2.0
    wire [11:0] v1047; shift_adder #(11, 11, 1, 1, 12, 0, 0) op_1047 (v219[10:0], v334[10:0], v1047[11:0]); // 2.0
    wire [12:0] v1048; shift_adder #(12, 12, 1, 1, 13, 0, 0) op_1048 (v389[11:0], v151[11:0], v1048[12:0]); // 2.0
    wire [10:0] v1049; shift_adder #(8, 11, 1, 1, 11, -1, 0) op_1049 (v65[7:0], v136[10:0], v1049[10:0]); // 2.0
    wire [25:0] v1050; shift_adder #(11, 11, 1, 1, 26, 15, 0) op_1050 (v155[10:0], v218[10:0], v1050[25:0]); // 2.0
    wire [32:0] v1051; shift_adder #(8, 16, 1, 1, 33, -24, 0) op_1051 (v106[7:0], v390[15:0], v1051[32:0]); // 2.0
    wire [14:0] v1052; shift_adder #(13, 9, 1, 1, 15, 5, 0) op_1052 (v391[12:0], v360[8:0], v1052[14:0]); // 2.0
    wire [14:0] v1053; shift_adder #(11, 12, 1, 1, 15, -4, 1) op_1053 (v294[10:0], v392[11:0], v1053[14:0]); // 2.0
    wire [10:0] v1054; shift_adder #(8, 11, 1, 1, 11, 0, 1) op_1054 (v65[7:0], v210[10:0], v1054[10:0]); // 2.0
    wire [14:0] v1055; shift_adder #(11, 11, 1, 1, 15, 4, 0) op_1055 (v200[10:0], v176[10:0], v1055[14:0]); // 2.0
    wire [11:0] v1056; shift_adder #(11, 10, 1, 1, 12, 1, 0) op_1056 (v352[10:0], v307[9:0], v1056[11:0]); // 2.0
    wire [13:0] v1057; shift_adder #(12, 14, 1, 1, 14, -1, 0) op_1057 (v279[11:0], v394[13:0], v1057[13:0]); // 2.0
    wire [23:0] v1058; shift_adder #(8, 11, 1, 1, 24, 13, 1) op_1058 (v85[7:0], v162[10:0], v1058[23:0]); // 2.0
    wire [18:0] v1059; shift_adder #(8, 10, 1, 1, 19, -10, 1) op_1059 (v72[7:0], v263[9:0], v1059[18:0]); // 2.0
    wire [32:0] v1060; shift_adder #(11, 11, 1, 1, 33, 22, 1) op_1060 (v386[10:0], v341[10:0], v1060[32:0]); // 2.0
    wire [21:0] v1061; shift_adder #(11, 16, 1, 1, 22, 6, 1) op_1061 (v283[10:0], v240[15:0], v1061[21:0]); // 2.0
    wire [20:0] v1062; shift_adder #(8, 12, 1, 1, 21, -12, 0) op_1062 (v100[7:0], v174[11:0], v1062[20:0]); // 2.0
    wire [16:0] v1063; shift_adder #(11, 11, 1, 1, 17, 6, 1) op_1063 (v132[10:0], v396[10:0], v1063[16:0]); // 2.0
    wire [15:0] v1064; shift_adder #(12, 12, 1, 1, 16, -4, 1) op_1064 (v397[11:0], v398[11:0], v1064[15:0]); // 2.0
    wire [34:0] v1065; shift_adder #(34, 17, 1, 1, 35, 18, 0) op_1065 (v399[33:0], v335[16:0], v1065[34:0]); // 2.0
    wire [14:0] v1066; shift_adder #(10, 11, 1, 1, 15, 4, 1) op_1066 (v307[9:0], v400[10:0], v1066[14:0]); // 2.0
    wire [21:0] v1067; shift_adder #(11, 20, 1, 1, 22, -11, 0) op_1067 (v300[10:0], v310[19:0], v1067[21:0]); // 2.0
    wire [11:0] v1068; shift_adder #(8, 11, 1, 1, 12, 1, 1) op_1068 (v111[7:0], v176[10:0], v1068[11:0]); // 2.0
    wire [11:0] v1069; shift_adder #(8, 11, 1, 1, 12, -2, 0) op_1069 (v102[7:0], v244[10:0], v1069[11:0]); // 2.0
    wire [12:0] v1070; shift_adder #(9, 12, 1, 1, 13, 1, 1) op_1070 (v401[8:0], v402[11:0], v1070[12:0]); // 2.0
    wire [14:0] v1071; shift_adder #(9, 11, 1, 1, 15, -5, 0) op_1071 (v403[8:0], v330[10:0], v1071[14:0]); // 2.0
    wire [13:0] v1072; shift_adder #(12, 12, 1, 1, 14, -2, 1) op_1072 (v292[11:0], v292[11:0], v1072[13:0]); // 2.0
    wire [17:0] v1073; shift_adder #(8, 11, 1, 1, 18, 7, 1) op_1073 (v72[7:0], v320[10:0], v1073[17:0]); // 2.0
    wire [12:0] v1074; shift_adder #(11, 11, 1, 1, 13, 2, 1) op_1074 (v218[10:0], v362[10:0], v1074[12:0]); // 2.0
    wire [19:0] v1075; shift_adder #(11, 11, 1, 1, 20, 9, 1) op_1075 (v228[10:0], v219[10:0], v1075[19:0]); // 2.0
    wire [25:0] v1076; shift_adder #(8, 11, 1, 1, 26, -17, 0) op_1076 (v79[7:0], v228[10:0], v1076[25:0]); // 2.0
    wire [11:0] v1077; shift_adder #(8, 11, 1, 1, 12, -2, 1) op_1077 (v120[7:0], v132[10:0], v1077[11:0]); // 2.0
    wire [12:0] v1078; shift_adder #(8, 11, 1, 1, 13, -4, 1) op_1078 (v75[7:0], v152[10:0], v1078[12:0]); // 2.0
    wire [12:0] v1079; shift_adder #(8, 11, 1, 1, 13, 2, 1) op_1079 (v103[7:0], v317[10:0], v1079[12:0]); // 2.0
    wire [11:0] v1080; shift_adder #(8, 11, 1, 1, 12, 1, 0) op_1080 (v101[7:0], v298[10:0], v1080[11:0]); // 2.0
    wire [10:0] v1081; shift_adder #(9, 9, 1, 1, 11, -1, 1) op_1081 (v322[8:0], v405[8:0], v1081[10:0]); // 2.0
    wire [11:0] v1082; shift_adder #(11, 11, 1, 1, 12, 0, 1) op_1082 (v163[10:0], v320[10:0], v1082[11:0]); // 2.0
    wire [12:0] v1083; shift_adder #(11, 12, 1, 1, 13, -1, 0) op_1083 (v312[10:0], v407[11:0], v1083[12:0]); // 2.0
    wire [14:0] v1084; shift_adder #(12, 12, 1, 1, 15, 3, 0) op_1084 (v204[11:0], v408[11:0], v1084[14:0]); // 2.0
    wire [13:0] v1085; shift_adder #(12, 12, 1, 1, 14, -2, 0) op_1085 (v321[11:0], v409[11:0], v1085[13:0]); // 2.0
    wire [12:0] v1086; shift_adder #(8, 13, 1, 1, 13, -2, 1) op_1086 (v70[7:0], v359[12:0], v1086[12:0]); // 2.0
    wire [23:0] v1087; shift_adder #(11, 12, 1, 1, 24, -13, 0) op_1087 (v245[10:0], v380[11:0], v1087[23:0]); // 2.0
    wire [15:0] v1088; shift_adder #(8, 11, 1, 1, 16, 5, 0) op_1088 (v127[7:0], v229[10:0], v1088[15:0]); // 2.0
    wire [15:0] v1089; shift_adder #(11, 11, 1, 1, 16, -5, 1) op_1089 (v156[10:0], v144[10:0], v1089[15:0]); // 2.0
    wire [20:0] v1090; shift_adder #(8, 11, 1, 1, 21, 10, 1) op_1090 (v109[7:0], v211[10:0], v1090[20:0]); // 2.0
    wire [15:0] v1091; shift_adder #(8, 14, 1, 1, 16, 2, 0) op_1091 (v84[7:0], v410[13:0], v1091[15:0]); // 2.0
    wire [24:0] v1092; shift_adder #(12, 12, 1, 1, 25, -13, 1) op_1092 (v174[11:0], v411[11:0], v1092[24:0]); // 2.0
    wire [29:0] v1093; shift_adder #(8, 14, 1, 1, 30, -21, 0) op_1093 (v101[7:0], v412[13:0], v1093[29:0]); // 2.0
    wire [17:0] v1094; shift_adder #(11, 11, 1, 1, 18, 7, 1) op_1094 (v134[10:0], v413[10:0], v1094[17:0]); // 2.0
    wire [24:0] v1095; shift_adder #(11, 17, 1, 1, 25, 8, 1) op_1095 (v210[10:0], v414[16:0], v1095[24:0]); // 2.0
    wire [17:0] v1096; shift_adder #(11, 12, 1, 1, 18, 6, 1) op_1096 (v134[10:0], v409[11:0], v1096[17:0]); // 2.0
    wire [12:0] v1097; shift_adder #(8, 11, 1, 1, 13, -4, 0) op_1097 (v105[7:0], v319[10:0], v1097[12:0]); // 2.0
    wire [15:0] v1098; shift_adder #(12, 11, 1, 1, 16, 5, 0) op_1098 (v151[11:0], v172[10:0], v1098[15:0]); // 2.0
    wire [17:0] v1099; shift_adder #(11, 11, 1, 1, 18, -7, 1) op_1099 (v229[10:0], v415[10:0], v1099[17:0]); // 2.0
    wire [11:0] v1100; shift_adder #(11, 11, 1, 1, 12, 0, 0) op_1100 (v181[10:0], v298[10:0], v1100[11:0]); // 2.0
    wire [19:0] v1101; shift_adder #(11, 11, 1, 1, 20, 9, 0) op_1101 (v142[10:0], v154[10:0], v1101[19:0]); // 2.0
    wire [11:0] v1102; shift_adder #(11, 12, 1, 1, 12, 0, 1) op_1102 (v185[10:0], v146[11:0], v1102[11:0]); // 2.0
    wire [11:0] v1103; shift_adder #(8, 11, 1, 1, 12, -2, 1) op_1103 (v98[7:0], v234[10:0], v1103[11:0]); // 2.0
    wire [13:0] v1104; shift_adder #(8, 11, 1, 1, 14, 3, 0) op_1104 (v94[7:0], v208[10:0], v1104[13:0]); // 2.0
    wire [11:0] v1105; shift_adder #(11, 11, 1, 1, 12, 1, 1) op_1105 (v338[10:0], v277[10:0], v1105[11:0]); // 2.0
    wire [15:0] v1106; shift_adder #(11, 12, 1, 1, 16, -5, 1) op_1106 (v386[10:0], v227[11:0], v1106[15:0]); // 2.0
    wire [14:0] v1107; shift_adder #(8, 12, 1, 1, 15, -6, 1) op_1107 (v89[7:0], v363[11:0], v1107[14:0]); // 2.0
    wire [14:0] v1108; shift_adder #(11, 13, 1, 1, 15, -4, 0) op_1108 (v139[10:0], v189[12:0], v1108[14:0]); // 2.0
    wire [14:0] v1109; shift_adder #(14, 11, 1, 1, 15, 3, 0) op_1109 (v417[13:0], v259[10:0], v1109[14:0]); // 2.0
    wire [33:0] v1110; shift_adder #(11, 11, 1, 1, 34, -23, 0) op_1110 (v134[10:0], v152[10:0], v1110[33:0]); // 2.0
    wire [13:0] v1111; shift_adder #(11, 13, 1, 1, 14, -2, 0) op_1111 (v276[10:0], v326[12:0], v1111[13:0]); // 2.0
    wire [13:0] v1112; shift_adder #(11, 13, 1, 1, 14, -2, 0) op_1112 (v139[10:0], v344[12:0], v1112[13:0]); // 2.0
    wire [18:0] v1113; shift_adder #(11, 10, 1, 1, 19, 9, 0) op_1113 (v232[10:0], v130[9:0], v1113[18:0]); // 2.0
    wire [15:0] v1114; shift_adder #(11, 11, 1, 1, 16, 5, 1) op_1114 (v131[10:0], v216[10:0], v1114[15:0]); // 2.0
    wire [10:0] v1115; shift_adder #(10, 11, 1, 1, 11, 0, 0) op_1115 (v419[9:0], v420[10:0], v1115[10:0]); // 2.0
    wire [13:0] v1116; shift_adder #(10, 14, 1, 1, 14, 0, 0) op_1116 (v421[9:0], v422[13:0], v1116[13:0]); // 2.0
    wire [13:0] v1117; shift_adder #(8, 9, 1, 1, 14, -5, 0) op_1117 (v126[7:0], v128[8:0], v1117[13:0]); // 2.0
    wire [16:0] v1118; shift_adder #(11, 11, 1, 1, 17, 6, 1) op_1118 (v228[10:0], v283[10:0], v1118[16:0]); // 2.0
    wire [14:0] v1119; shift_adder #(8, 11, 1, 1, 15, -6, 0) op_1119 (v119[7:0], v181[10:0], v1119[14:0]); // 2.0
    wire [14:0] v1120; shift_adder #(8, 12, 1, 1, 15, -6, 0) op_1120 (v113[7:0], v423[11:0], v1120[14:0]); // 2.0
    wire [11:0] v1121; shift_adder #(8, 11, 1, 1, 12, -3, 1) op_1121 (v107[7:0], v379[10:0], v1121[11:0]); // 2.0
    wire [10:0] v1122; shift_adder #(8, 11, 1, 1, 11, -1, 1) op_1122 (v64[7:0], v229[10:0], v1122[10:0]); // 2.0
    wire [12:0] v1123; shift_adder #(11, 11, 1, 1, 13, 2, 0) op_1123 (v424[10:0], v425[10:0], v1123[12:0]); // 2.0
    wire [14:0] v1124; shift_adder #(8, 11, 1, 1, 15, 4, 0) op_1124 (v82[7:0], v173[10:0], v1124[14:0]); // 2.0
    wire [11:0] v1125; shift_adder #(11, 11, 1, 1, 12, 1, 0) op_1125 (v217[10:0], v418[10:0], v1125[11:0]); // 2.0
    wire [13:0] v1126; shift_adder #(8, 11, 1, 1, 14, 3, 1) op_1126 (v116[7:0], v289[10:0], v1126[13:0]); // 2.0
    wire [14:0] v1127; shift_adder #(11, 11, 1, 1, 15, -4, 1) op_1127 (v264[10:0], v181[10:0], v1127[14:0]); // 2.0
    wire [20:0] v1128; shift_adder #(11, 11, 1, 1, 21, -10, 1) op_1128 (v338[10:0], v320[10:0], v1128[20:0]); // 2.0
    wire [14:0] v1129; shift_adder #(14, 11, 1, 1, 15, 4, 0) op_1129 (v417[13:0], v274[10:0], v1129[14:0]); // 2.0
    wire [17:0] v1130; shift_adder #(8, 12, 1, 1, 18, 6, 1) op_1130 (v71[7:0], v239[11:0], v1130[17:0]); // 2.0
    wire [22:0] v1131; shift_adder #(11, 11, 1, 1, 23, -12, 1) op_1131 (v229[10:0], v259[10:0], v1131[22:0]); // 2.0
    wire [13:0] v1132; shift_adder #(11, 11, 1, 1, 14, -3, 1) op_1132 (v140[10:0], v293[10:0], v1132[13:0]); // 2.0
    wire [21:0] v1133; shift_adder #(21, 13, 1, 1, 22, 9, 0) op_1133 (v427[20:0], v359[12:0], v1133[21:0]); // 2.0
    wire [12:0] v1134; shift_adder #(11, 12, 1, 1, 13, -2, 1) op_1134 (v145[10:0], v365[11:0], v1134[12:0]); // 2.0
    wire [13:0] v1135; shift_adder #(8, 11, 1, 1, 14, 3, 1) op_1135 (v114[7:0], v228[10:0], v1135[13:0]); // 2.0
    wire [11:0] v1136; shift_adder #(11, 11, 1, 1, 12, 1, 0) op_1136 (v223[10:0], v200[10:0], v1136[11:0]); // 2.0
    wire [10:0] v1137; shift_adder #(8, 10, 1, 1, 11, 1, 0) op_1137 (v95[7:0], v428[9:0], v1137[10:0]); // 2.0
    wire [12:0] v1138; shift_adder #(8, 12, 1, 1, 13, 1, 1) op_1138 (v124[7:0], v247[11:0], v1138[12:0]); // 2.0
    wire [13:0] v1139; shift_adder #(8, 11, 1, 1, 14, -5, 1) op_1139 (v124[7:0], v139[10:0], v1139[13:0]); // 2.0
    wire [30:0] v1140; shift_adder #(11, 11, 1, 1, 31, 20, 1) op_1140 (v358[10:0], v187[10:0], v1140[30:0]); // 2.0
    wire [22:0] v1141; shift_adder #(8, 11, 1, 1, 23, -14, 0) op_1141 (v113[7:0], v289[10:0], v1141[22:0]); // 2.0
    wire [19:0] v1142; shift_adder #(11, 12, 1, 1, 20, -9, 0) op_1142 (v245[10:0], v202[11:0], v1142[19:0]); // 2.0
    wire [18:0] v1143; shift_adder #(18, 11, 1, 1, 19, 8, 0) op_1143 (v429[17:0], v320[10:0], v1143[18:0]); // 2.0
    wire [20:0] v1144; shift_adder #(11, 11, 1, 1, 21, -10, 1) op_1144 (v147[10:0], v430[10:0], v1144[20:0]); // 2.0
    wire [30:0] v1145; shift_adder #(8, 10, 1, 1, 31, -22, 1) op_1145 (v105[7:0], v254[9:0], v1145[30:0]); // 2.0
    wire [16:0] v1146; shift_adder #(8, 11, 1, 1, 17, 6, 0) op_1146 (v116[7:0], v132[10:0], v1146[16:0]); // 2.0
    wire [11:0] v1147; shift_adder #(11, 11, 1, 1, 12, 0, 1) op_1147 (v216[10:0], v163[10:0], v1147[11:0]); // 2.0
    wire [20:0] v1148; shift_adder #(19, 10, 1, 1, 21, 11, 0) op_1148 (v315[18:0], v432[9:0], v1148[20:0]); // 2.0
    wire [23:0] v1149; shift_adder #(11, 9, 1, 1, 24, 14, 0) op_1149 (v362[10:0], v433[8:0], v1149[23:0]); // 2.0
    wire [17:0] v1150; shift_adder #(12, 12, 1, 1, 18, -6, 1) op_1150 (v434[11:0], v314[11:0], v1150[17:0]); // 2.0
    wire [16:0] v1151; shift_adder #(11, 11, 1, 1, 17, 6, 0) op_1151 (v158[10:0], v270[10:0], v1151[16:0]); // 2.0
    wire [15:0] v1152; shift_adder #(11, 12, 1, 1, 16, 4, 0) op_1152 (v216[10:0], v174[11:0], v1152[15:0]); // 2.0
    wire [11:0] v1153; shift_adder #(11, 11, 1, 1, 12, -1, 0) op_1153 (v362[10:0], v420[10:0], v1153[11:0]); // 2.0
    wire [16:0] v1154; shift_adder #(12, 10, 1, 1, 17, 7, 1) op_1154 (v292[11:0], v282[9:0], v1154[16:0]); // 2.0
    wire [11:0] v1155; shift_adder #(11, 11, 1, 1, 12, 0, 0) op_1155 (v228[10:0], v171[10:0], v1155[11:0]); // 2.0
    wire [15:0] v1156; shift_adder #(11, 11, 1, 1, 16, -5, 1) op_1156 (v144[10:0], v362[10:0], v1156[15:0]); // 2.0
    wire [16:0] v1157; shift_adder #(10, 17, 1, 1, 17, 0, 1) op_1157 (v435[9:0], v436[16:0], v1157[16:0]); // 2.0
    wire [14:0] v1158; shift_adder #(12, 10, 1, 1, 15, 5, 0) op_1158 (v292[11:0], v437[9:0], v1158[14:0]); // 2.0
    wire [11:0] v1159; shift_adder #(11, 11, 1, 1, 12, -1, 0) op_1159 (v179[10:0], v301[10:0], v1159[11:0]); // 2.0
    wire [11:0] v1160; shift_adder #(8, 11, 1, 1, 12, -3, 0) op_1160 (v80[7:0], v171[10:0], v1160[11:0]); // 2.0
    wire [10:0] v1161; shift_adder #(8, 11, 1, 1, 11, 0, 1) op_1161 (v104[7:0], v162[10:0], v1161[10:0]); // 2.0
    wire [13:0] v1162; shift_adder #(11, 11, 1, 1, 14, 3, 0) op_1162 (v237[10:0], v210[10:0], v1162[13:0]); // 2.0
    wire [12:0] v1163; shift_adder #(11, 12, 1, 1, 13, -1, 1) op_1163 (v270[10:0], v438[11:0], v1163[12:0]); // 2.0
    wire [12:0] v1164; shift_adder #(13, 11, 1, 1, 13, 1, 0) op_1164 (v192[12:0], v150[10:0], v1164[12:0]); // 2.0
    wire [13:0] v1165; shift_adder #(8, 11, 1, 1, 14, 3, 0) op_1165 (v124[7:0], v374[10:0], v1165[13:0]); // 2.0
    wire [28:0] v1166; shift_adder #(12, 29, 1, 1, 29, -2, 1) op_1166 (v387[11:0], v439[28:0], v1166[28:0]); // 2.0
    wire [25:0] v1167; shift_adder #(11, 11, 1, 1, 26, 15, 1) op_1167 (v206[10:0], v277[10:0], v1167[25:0]); // 2.0
    wire [20:0] v1168; shift_adder #(8, 11, 1, 1, 21, -12, 0) op_1168 (v127[7:0], v132[10:0], v1168[20:0]); // 2.0
    wire [15:0] v1169; shift_adder #(11, 12, 1, 1, 16, -5, 1) op_1169 (v211[10:0], v387[11:0], v1169[15:0]); // 2.0
    wire [11:0] v1170; shift_adder #(11, 11, 1, 1, 12, -1, 0) op_1170 (v141[10:0], v358[10:0], v1170[11:0]); // 2.0
    wire [11:0] v1171; shift_adder #(11, 11, 1, 1, 12, 0, 1) op_1171 (v317[10:0], v173[10:0], v1171[11:0]); // 2.0
    wire [23:0] v1172; shift_adder #(23, 12, 1, 1, 24, 11, 0) op_1172 (v440[22:0], v355[11:0], v1172[23:0]); // 2.0
    wire [14:0] v1173; shift_adder #(11, 12, 1, 1, 15, -4, 1) op_1173 (v190[10:0], v383[11:0], v1173[14:0]); // 2.0
    wire [10:0] v1174; shift_adder #(9, 10, 1, 1, 11, -1, 0) op_1174 (v441[8:0], v442[9:0], v1174[10:0]); // 2.0
    wire [16:0] v1175; shift_adder #(11, 11, 1, 1, 17, 6, 0) op_1175 (v232[10:0], v212[10:0], v1175[16:0]); // 2.0
    wire [11:0] v1176; shift_adder #(11, 11, 1, 1, 12, 0, 0) op_1176 (v246[10:0], v443[10:0], v1176[11:0]); // 2.0
    wire [12:0] v1177; shift_adder #(11, 11, 1, 1, 13, 2, 0) op_1177 (v191[10:0], v425[10:0], v1177[12:0]); // 2.0
    wire [11:0] v1178; shift_adder #(8, 11, 1, 1, 12, 1, 1) op_1178 (v73[7:0], v266[10:0], v1178[11:0]); // 2.0
    wire [21:0] v1179; shift_adder #(8, 11, 1, 1, 22, 11, 1) op_1179 (v74[7:0], v283[10:0], v1179[21:0]); // 2.0
    wire [12:0] v1180; shift_adder #(11, 11, 1, 1, 13, -2, 1) op_1180 (v171[10:0], v319[10:0], v1180[12:0]); // 2.0
    wire [20:0] v1181; shift_adder #(11, 11, 1, 1, 21, -10, 0) op_1181 (v338[10:0], v165[10:0], v1181[20:0]); // 2.0
    wire [11:0] v1182; shift_adder #(11, 11, 1, 1, 12, -1, 0) op_1182 (v168[10:0], v420[10:0], v1182[11:0]); // 2.0
    wire [14:0] v1183; shift_adder #(11, 14, 1, 1, 15, -3, 0) op_1183 (v353[10:0], v444[13:0], v1183[14:0]); // 2.0
    wire [12:0] v1184; shift_adder #(12, 10, 1, 1, 13, 2, 0) op_1184 (v305[11:0], v445[9:0], v1184[12:0]); // 2.0
    wire [10:0] v1185; shift_adder #(10, 9, 1, 1, 11, 1, 0) op_1185 (v291[9:0], v401[8:0], v1185[10:0]); // 2.0
    wire [14:0] v1186; shift_adder #(8, 11, 1, 1, 15, 4, 1) op_1186 (v81[7:0], v361[10:0], v1186[14:0]); // 2.0
    wire [12:0] v1187; shift_adder #(8, 12, 1, 1, 13, -3, 0) op_1187 (v118[7:0], v314[11:0], v1187[12:0]); // 2.0
    wire [11:0] v1188; shift_adder #(11, 11, 1, 1, 12, 0, 1) op_1188 (v173[10:0], v182[10:0], v1188[11:0]); // 2.0
    wire [12:0] v1189; shift_adder #(8, 11, 1, 1, 13, 2, 1) op_1189 (v80[7:0], v144[10:0], v1189[12:0]); // 2.0
    wire [11:0] v1190; shift_adder #(11, 11, 1, 1, 12, -1, 1) op_1190 (v136[10:0], v168[10:0], v1190[11:0]); // 2.0
    wire [20:0] v1191; shift_adder #(8, 11, 1, 1, 21, -12, 1) op_1191 (v64[7:0], v148[10:0], v1191[20:0]); // 2.0
    wire [21:0] v1192; shift_adder #(11, 9, 1, 1, 22, -11, 0) op_1192 (v275[10:0], v221[8:0], v1192[21:0]); // 2.0
    wire [31:0] v1193; shift_adder #(32, 11, 1, 1, 32, 17, 0) op_1193 (v448[31:0], v135[10:0], v1193[31:0]); // 2.0
    wire [24:0] v1194; shift_adder #(11, 11, 1, 1, 25, -14, 1) op_1194 (v158[10:0], v255[10:0], v1194[24:0]); // 2.0
    wire [18:0] v1195; shift_adder #(8, 11, 1, 1, 19, 8, 1) op_1195 (v115[7:0], v211[10:0], v1195[18:0]); // 2.0
    wire [11:0] v1196; shift_adder #(11, 11, 1, 1, 12, -1, 0) op_1196 (v148[10:0], v154[10:0], v1196[11:0]); // 2.0
    wire [20:0] v1197; shift_adder #(11, 11, 1, 1, 21, -10, 0) op_1197 (v362[10:0], v142[10:0], v1197[20:0]); // 2.0
    wire [18:0] v1198; shift_adder #(8, 10, 1, 1, 19, -10, 0) op_1198 (v98[7:0], v450[9:0], v1198[18:0]); // 2.0
    wire [11:0] v1199; shift_adder #(8, 11, 1, 1, 12, -3, 0) op_1199 (v99[7:0], v193[10:0], v1199[11:0]); // 2.0
    wire [22:0] v1200; shift_adder #(8, 13, 1, 1, 23, 10, 1) op_1200 (v97[7:0], v451[12:0], v1200[22:0]); // 2.0
    wire [15:0] v1201; shift_adder #(11, 12, 1, 1, 16, -5, 0) op_1201 (v144[10:0], v372[11:0], v1201[15:0]); // 2.0
    wire [12:0] v1202; shift_adder #(11, 11, 1, 1, 13, 2, 1) op_1202 (v155[10:0], v175[10:0], v1202[12:0]); // 2.0
    wire [11:0] v1203; shift_adder #(11, 11, 1, 1, 12, 1, 0) op_1203 (v312[10:0], v393[10:0], v1203[11:0]); // 2.0
    wire [13:0] v1204; shift_adder #(12, 11, 1, 1, 14, -2, 0) op_1204 (v452[11:0], v195[10:0], v1204[13:0]); // 2.0
    wire [14:0] v1205; shift_adder #(11, 11, 1, 1, 15, 4, 1) op_1205 (v238[10:0], v133[10:0], v1205[14:0]); // 2.0
    wire [20:0] v1206; shift_adder #(14, 21, 1, 1, 21, -4, 0) op_1206 (v454[13:0], v427[20:0], v1206[20:0]); // 2.0
    wire [17:0] v1207; shift_adder #(15, 11, 1, 1, 18, 7, 0) op_1207 (v456[14:0], v215[10:0], v1207[17:0]); // 2.0
    wire [17:0] v1208; shift_adder #(11, 12, 1, 1, 18, -7, 1) op_1208 (v375[10:0], v457[11:0], v1208[17:0]); // 2.0
    wire [12:0] v1209; shift_adder #(11, 12, 1, 1, 13, -1, 1) op_1209 (v234[10:0], v387[11:0], v1209[12:0]); // 2.0
    wire [18:0] v1210; shift_adder #(8, 19, 1, 1, 19, 0, 0) op_1210 (v126[7:0], v376[18:0], v1210[18:0]); // 2.0
    wire [11:0] v1211; shift_adder #(11, 11, 1, 1, 12, 0, 0) op_1211 (v241[10:0], v353[10:0], v1211[11:0]); // 2.0
    wire [20:0] v1212; shift_adder #(11, 12, 1, 1, 21, 9, 0) op_1212 (v148[10:0], v438[11:0], v1212[20:0]); // 2.0
    wire [15:0] v1213; shift_adder #(8, 11, 1, 1, 16, 5, 0) op_1213 (v105[7:0], v195[10:0], v1213[15:0]); // 2.0
    wire [11:0] v1214; shift_adder #(11, 11, 1, 1, 12, 1, 0) op_1214 (v203[10:0], v215[10:0], v1214[11:0]); // 2.0
    wire [22:0] v1215; shift_adder #(11, 13, 1, 1, 23, -12, 1) op_1215 (v232[10:0], v458[12:0], v1215[22:0]); // 2.0
    wire [20:0] v1216; shift_adder #(8, 10, 1, 1, 21, 11, 0) op_1216 (v69[7:0], v459[9:0], v1216[20:0]); // 2.0
    wire [18:0] v1217; shift_adder #(8, 11, 1, 1, 19, -10, 0) op_1217 (v127[7:0], v148[10:0], v1217[18:0]); // 2.0
    wire [18:0] v1218; shift_adder #(11, 14, 1, 1, 19, 5, 1) op_1218 (v155[10:0], v460[13:0], v1218[18:0]); // 2.0
    wire [28:0] v1219; shift_adder #(8, 9, 1, 1, 29, 19, 1) op_1219 (v109[7:0], v395[8:0], v1219[28:0]); // 2.0
    wire [16:0] v1220; shift_adder #(11, 11, 1, 1, 17, 6, 1) op_1220 (v219[10:0], v200[10:0], v1220[16:0]); // 2.0
    wire [16:0] v1221; shift_adder #(8, 10, 1, 1, 17, -8, 0) op_1221 (v106[7:0], v366[9:0], v1221[16:0]); // 2.0
    wire [13:0] v1222; shift_adder #(8, 11, 1, 1, 14, -5, 1) op_1222 (v66[7:0], v136[10:0], v1222[13:0]); // 2.0
    wire [29:0] v1223; shift_adder #(11, 11, 1, 1, 30, 19, 1) op_1223 (v228[10:0], v155[10:0], v1223[29:0]); // 2.0
    wire [19:0] v1224; shift_adder #(11, 11, 1, 1, 20, 9, 1) op_1224 (v298[10:0], v191[10:0], v1224[19:0]); // 2.0
    wire [14:0] v1225; shift_adder #(12, 14, 1, 1, 15, 1, 0) op_1225 (v184[11:0], v454[13:0], v1225[14:0]); // 2.0
    wire [18:0] v1226; shift_adder #(11, 12, 1, 1, 19, 7, 1) op_1226 (v246[10:0], v333[11:0], v1226[18:0]); // 2.0
    wire [12:0] v1227; shift_adder #(8, 11, 1, 1, 13, -4, 0) op_1227 (v78[7:0], v294[10:0], v1227[12:0]); // 2.0
    wire [13:0] v1228; shift_adder #(11, 9, 1, 1, 14, 4, 0) op_1228 (v362[10:0], v231[8:0], v1228[13:0]); // 2.0
    wire [13:0] v1229; shift_adder #(8, 11, 1, 1, 14, 3, 0) op_1229 (v97[7:0], v312[10:0], v1229[13:0]); // 2.0
    wire [12:0] v1230; shift_adder #(11, 12, 1, 1, 13, 1, 1) op_1230 (v420[10:0], v382[11:0], v1230[12:0]); // 2.0
    wire [16:0] v1231; shift_adder #(8, 11, 1, 1, 17, 6, 0) op_1231 (v125[7:0], v182[10:0], v1231[16:0]); // 2.0
    wire [29:0] v1232; shift_adder #(12, 12, 1, 1, 30, 18, 0) op_1232 (v333[11:0], v288[11:0], v1232[29:0]); // 2.0
    wire [13:0] v1233; shift_adder #(12, 10, 1, 1, 14, 3, 0) op_1233 (v462[11:0], v463[9:0], v1233[13:0]); // 2.0
    wire [11:0] v1234; shift_adder #(8, 12, 1, 1, 12, -1, 1) op_1234 (v116[7:0], v464[11:0], v1234[11:0]); // 2.0
    wire [17:0] v1235; shift_adder #(8, 11, 1, 1, 18, -9, 1) op_1235 (v73[7:0], v168[10:0], v1235[17:0]); // 2.0
    wire [16:0] v1236; shift_adder #(8, 15, 1, 1, 17, -8, 0) op_1236 (v121[7:0], v465[14:0], v1236[16:0]); // 2.0
    wire [18:0] v1237; shift_adder #(12, 18, 1, 1, 19, -6, 1) op_1237 (v243[11:0], v286[17:0], v1237[18:0]); // 2.0
    wire [15:0] v1238; shift_adder #(8, 11, 1, 1, 16, 5, 0) op_1238 (v72[7:0], v158[10:0], v1238[15:0]); // 2.0
    wire [29:0] v1239; shift_adder #(11, 13, 1, 1, 30, 17, 1) op_1239 (v455[10:0], v149[12:0], v1239[29:0]); // 2.0
    wire [10:0] v1240; shift_adder #(10, 9, 1, 1, 11, 0, 0) op_1240 (v466[9:0], v467[8:0], v1240[10:0]); // 2.0
    wire [11:0] v1241; shift_adder #(10, 11, 1, 1, 12, 1, 0) op_1241 (v468[9:0], v215[10:0], v1241[11:0]); // 2.0
    wire [11:0] v1242; shift_adder #(10, 11, 1, 1, 12, -1, 0) op_1242 (v469[9:0], v168[10:0], v1242[11:0]); // 2.0
    wire [27:0] v1243; shift_adder #(11, 12, 1, 1, 28, 16, 1) op_1243 (v188[10:0], v333[11:0], v1243[27:0]); // 2.0
    wire [11:0] v1244; shift_adder #(11, 11, 1, 1, 12, 1, 0) op_1244 (v188[10:0], v178[10:0], v1244[11:0]); // 2.0
    wire [27:0] v1245; shift_adder #(11, 11, 1, 1, 28, 17, 0) op_1245 (v182[10:0], v191[10:0], v1245[27:0]); // 2.0
    wire [26:0] v1246; shift_adder #(11, 10, 1, 1, 27, 17, 1) op_1246 (v396[10:0], v130[9:0], v1246[26:0]); // 2.0
    wire [12:0] v1247; shift_adder #(8, 12, 1, 1, 13, -3, 1) op_1247 (v101[7:0], v473[11:0], v1247[12:0]); // 2.0
    wire [14:0] v1248; shift_adder #(9, 14, 1, 1, 15, -5, 0) op_1248 (v360[8:0], v474[13:0], v1248[14:0]); // 2.0
    wire [15:0] v1249; shift_adder #(11, 16, 1, 1, 16, -3, 1) op_1249 (v244[10:0], v166[15:0], v1249[15:0]); // 2.0
    wire [13:0] v1250; shift_adder #(11, 12, 1, 1, 14, 2, 1) op_1250 (v147[10:0], v174[11:0], v1250[13:0]); // 2.0
    wire [13:0] v1251; shift_adder #(12, 13, 1, 1, 14, -2, 0) op_1251 (v475[11:0], v476[12:0], v1251[13:0]); // 2.0
    wire [14:0] v1252; shift_adder #(11, 11, 1, 1, 15, -4, 0) op_1252 (v150[10:0], v150[10:0], v1252[14:0]); // 2.0
    wire [11:0] v1253; shift_adder #(11, 11, 1, 1, 12, 0, 0) op_1253 (v218[10:0], v157[10:0], v1253[11:0]); // 2.0
    wire [14:0] v1254; shift_adder #(11, 11, 1, 1, 15, -4, 0) op_1254 (v200[10:0], v328[10:0], v1254[14:0]); // 2.0
    wire [11:0] v1255; shift_adder #(11, 11, 1, 1, 12, 0, 1) op_1255 (v190[10:0], v139[10:0], v1255[11:0]); // 2.0
    wire [13:0] v1256; shift_adder #(11, 10, 1, 1, 14, 4, 0) op_1256 (v190[10:0], v248[9:0], v1256[13:0]); // 2.0
    wire [11:0] v1257; shift_adder #(9, 11, 1, 1, 12, -1, 0) op_1257 (v477[8:0], v478[10:0], v1257[11:0]); // 2.0
    wire [11:0] v1258; shift_adder #(9, 11, 1, 1, 12, -2, 0) op_1258 (v479[8:0], v217[10:0], v1258[11:0]); // 2.0
    wire [11:0] v1259; shift_adder #(11, 11, 1, 1, 12, 0, 0) op_1259 (v317[10:0], v181[10:0], v1259[11:0]); // 2.0
    wire [26:0] v1260; shift_adder #(8, 27, 1, 1, 27, -17, 1) op_1260 (v108[7:0], v480[26:0], v1260[26:0]); // 2.0
    wire [11:0] v1261; shift_adder #(8, 11, 1, 1, 12, -3, 1) op_1261 (v112[7:0], v133[10:0], v1261[11:0]); // 2.0
    wire [11:0] v1262; shift_adder #(8, 11, 1, 1, 12, -3, 0) op_1262 (v125[7:0], v289[10:0], v1262[11:0]); // 2.0
    wire [12:0] v1263; shift_adder #(11, 11, 1, 1, 13, -2, 1) op_1263 (v297[10:0], v153[10:0], v1263[12:0]); // 2.0
    wire [23:0] v1264; shift_adder #(11, 11, 1, 1, 24, 13, 1) op_1264 (v228[10:0], v223[10:0], v1264[23:0]); // 2.0
    wire [14:0] v1265; shift_adder #(8, 11, 1, 1, 15, 4, 0) op_1265 (v110[7:0], v297[10:0], v1265[14:0]); // 2.0
    wire [20:0] v1266; shift_adder #(11, 11, 1, 1, 21, 10, 1) op_1266 (v245[10:0], v145[10:0], v1266[20:0]); // 2.0
    wire [20:0] v1267; shift_adder #(14, 15, 1, 1, 21, -7, 0) op_1267 (v481[13:0], v482[14:0], v1267[20:0]); // 2.0
    wire [23:0] v1268; shift_adder #(11, 11, 1, 1, 24, 13, 1) op_1268 (v206[10:0], v161[10:0], v1268[23:0]); // 2.0
    wire [24:0] v1269; shift_adder #(11, 12, 1, 1, 25, -14, 1) op_1269 (v155[10:0], v305[11:0], v1269[24:0]); // 2.0
    wire [13:0] v1270; shift_adder #(11, 11, 1, 1, 14, -3, 0) op_1270 (v141[10:0], v294[10:0], v1270[13:0]); // 2.0
    wire [26:0] v1271; shift_adder #(11, 14, 1, 1, 27, 13, 1) op_1271 (v216[10:0], v483[13:0], v1271[26:0]); // 2.0
    wire [14:0] v1272; shift_adder #(11, 11, 1, 1, 15, 4, 1) op_1272 (v276[10:0], v131[10:0], v1272[14:0]); // 2.0
    wire [10:0] v1273; shift_adder #(8, 11, 1, 1, 11, 0, 1) op_1273 (v67[7:0], v188[10:0], v1273[10:0]); // 2.0
    wire [26:0] v1274; shift_adder #(11, 12, 1, 1, 27, -16, 1) op_1274 (v244[10:0], v409[11:0], v1274[26:0]); // 2.0
    wire [15:0] v1275; shift_adder #(11, 11, 1, 1, 16, -5, 0) op_1275 (v275[10:0], v259[10:0], v1275[15:0]); // 2.0
    wire [11:0] v1276; shift_adder #(8, 11, 1, 1, 12, -3, 1) op_1276 (v120[7:0], v210[10:0], v1276[11:0]); // 2.0
    wire [11:0] v1277; shift_adder #(11, 11, 1, 1, 12, -1, 1) op_1277 (v182[10:0], v329[10:0], v1277[11:0]); // 2.0
    wire [11:0] v1278; shift_adder #(11, 11, 1, 1, 12, -1, 1) op_1278 (v277[10:0], v165[10:0], v1278[11:0]); // 2.0
    wire [12:0] v1279; shift_adder #(8, 11, 1, 1, 13, 2, 1) op_1279 (v115[7:0], v283[10:0], v1279[12:0]); // 2.0
    wire [12:0] v1280; shift_adder #(8, 11, 1, 1, 13, -4, 0) op_1280 (v95[7:0], v425[10:0], v1280[12:0]); // 2.0
    wire [13:0] v1281; shift_adder #(8, 11, 1, 1, 14, 3, 0) op_1281 (v121[7:0], v132[10:0], v1281[13:0]); // 2.0
    wire [14:0] v1282; shift_adder #(11, 11, 1, 1, 15, -4, 0) op_1282 (v163[10:0], v418[10:0], v1282[14:0]); // 2.0
    wire [11:0] v1283; shift_adder #(8, 11, 1, 1, 12, 1, 1) op_1283 (v66[7:0], v169[10:0], v1283[11:0]); // 2.0
    wire [10:0] v1284; shift_adder #(8, 11, 1, 1, 11, -1, 0) op_1284 (v108[7:0], v177[10:0], v1284[10:0]); // 2.0
    wire [14:0] v1285; shift_adder #(11, 11, 1, 1, 15, -4, 0) op_1285 (v199[10:0], v199[10:0], v1285[14:0]); // 2.0
    wire [19:0] v1286; shift_adder #(11, 11, 1, 1, 20, 9, 0) op_1286 (v229[10:0], v185[10:0], v1286[19:0]); // 2.0
    wire [23:0] v1287; shift_adder #(11, 11, 1, 1, 24, -13, 1) op_1287 (v173[10:0], v367[10:0], v1287[23:0]); // 2.0
    wire [13:0] v1288; shift_adder #(11, 11, 1, 1, 14, -3, 1) op_1288 (v237[10:0], v244[10:0], v1288[13:0]); // 2.0
    wire [19:0] v1289; shift_adder #(8, 11, 1, 1, 20, 9, 1) op_1289 (v122[7:0], v144[10:0], v1289[19:0]); // 2.0
    wire [13:0] v1290; shift_adder #(11, 12, 1, 1, 14, -3, 0) op_1290 (v140[10:0], v473[11:0], v1290[13:0]); // 2.0
    wire [16:0] v1291; shift_adder #(8, 11, 1, 1, 17, 6, 0) op_1291 (v99[7:0], v301[10:0], v1291[16:0]); // 2.0
    wire [18:0] v1292; shift_adder #(19, 10, 1, 1, 19, 8, 0) op_1292 (v485[18:0], v428[9:0], v1292[18:0]); // 2.0
    wire [10:0] v1293; shift_adder #(11, 10, 1, 1, 11, 0, 0) op_1293 (v216[10:0], v260[9:0], v1293[10:0]); // 2.0
    wire [12:0] v1294; shift_adder #(9, 11, 1, 1, 13, -3, 0) op_1294 (v486[8:0], v487[10:0], v1294[12:0]); // 2.0
    wire [12:0] v1295; shift_adder #(11, 11, 1, 1, 13, 2, 0) op_1295 (v141[10:0], v276[10:0], v1295[12:0]); // 2.0
    wire [14:0] v1296; shift_adder #(14, 11, 1, 1, 15, 3, 0) op_1296 (v488[13:0], v191[10:0], v1296[14:0]); // 2.0
    wire [22:0] v1297; shift_adder #(8, 12, 1, 1, 23, 11, 0) op_1297 (v103[7:0], v305[11:0], v1297[22:0]); // 2.0
    wire [10:0] v1298; shift_adder #(11, 10, 1, 1, 11, 0, 1) op_1298 (v245[10:0], v225[9:0], v1298[10:0]); // 2.0
    wire [13:0] v1299; shift_adder #(11, 11, 1, 1, 14, -3, 1) op_1299 (v206[10:0], v268[10:0], v1299[13:0]); // 2.0
    wire [13:0] v1300; shift_adder #(11, 11, 1, 1, 14, 3, 0) op_1300 (v250[10:0], v242[10:0], v1300[13:0]); // 2.0
    wire [13:0] v1301; shift_adder #(11, 12, 1, 1, 14, 2, 1) op_1301 (v362[10:0], v243[11:0], v1301[13:0]); // 2.0
    wire [19:0] v1302; shift_adder #(11, 11, 1, 1, 20, -9, 0) op_1302 (v386[10:0], v242[10:0], v1302[19:0]); // 2.0
    wire [13:0] v1303; shift_adder #(8, 9, 1, 1, 14, 4, 0) op_1303 (v122[7:0], v351[8:0], v1303[13:0]); // 2.0
    wire [14:0] v1304; shift_adder #(8, 14, 1, 1, 15, 1, 1) op_1304 (v67[7:0], v472[13:0], v1304[14:0]); // 2.0
    wire [11:0] v1305; shift_adder #(9, 11, 1, 1, 12, -2, 0) op_1305 (v309[8:0], v275[10:0], v1305[11:0]); // 2.0
    wire [10:0] v1306; shift_adder #(8, 11, 1, 1, 11, -1, 1) op_1306 (v70[7:0], v211[10:0], v1306[10:0]); // 2.0
    wire [13:0] v1307; shift_adder #(11, 11, 1, 1, 14, -3, 1) op_1307 (v199[10:0], v430[10:0], v1307[13:0]); // 2.0
    wire [11:0] v1308; shift_adder #(11, 11, 1, 1, 12, 0, 0) op_1308 (v201[10:0], v377[10:0], v1308[11:0]); // 2.0
    wire [11:0] v1309; shift_adder #(11, 11, 1, 1, 12, 0, 0) op_1309 (v237[10:0], v294[10:0], v1309[11:0]); // 2.0
    wire [13:0] v1310; shift_adder #(11, 10, 1, 1, 14, 4, 0) op_1310 (v242[10:0], v489[9:0], v1310[13:0]); // 2.0
    wire [15:0] v1311; shift_adder #(8, 13, 1, 1, 16, -7, 0) op_1311 (v122[7:0], v149[12:0], v1311[15:0]); // 2.0
    wire [16:0] v1312; shift_adder #(8, 9, 1, 1, 17, -8, 1) op_1312 (v114[7:0], v138[8:0], v1312[16:0]); // 2.0
    wire [13:0] v1313; shift_adder #(11, 11, 1, 1, 14, 3, 1) op_1313 (v155[10:0], v216[10:0], v1313[13:0]); // 2.0
    wire [11:0] v1314; shift_adder #(12, 11, 1, 1, 12, 0, 0) op_1314 (v411[11:0], v491[10:0], v1314[11:0]); // 2.0
    wire [16:0] v1315; shift_adder #(11, 11, 1, 1, 17, 6, 1) op_1315 (v418[10:0], v424[10:0], v1315[16:0]); // 2.0
    wire [17:0] v1316; shift_adder #(11, 11, 1, 1, 18, 7, 0) op_1316 (v156[10:0], v234[10:0], v1316[17:0]); // 2.0
    wire [13:0] v1317; shift_adder #(8, 12, 1, 1, 14, 2, 1) op_1317 (v103[7:0], v151[11:0], v1317[13:0]); // 2.0
    wire [31:0] v1318; shift_adder #(8, 11, 1, 1, 32, 21, 1) op_1318 (v123[7:0], v338[10:0], v1318[31:0]); // 2.0
    wire [22:0] v1319; shift_adder #(11, 11, 1, 1, 23, 12, 0) op_1319 (v133[10:0], v176[10:0], v1319[22:0]); // 2.0
    wire [18:0] v1320; shift_adder #(11, 11, 1, 1, 19, -8, 1) op_1320 (v328[10:0], v328[10:0], v1320[18:0]); // 2.0
    wire [18:0] v1321; shift_adder #(11, 11, 1, 1, 19, -8, 1) op_1321 (v172[10:0], v232[10:0], v1321[18:0]); // 2.0
    wire [32:0] v1322; shift_adder #(11, 11, 1, 1, 33, 22, 0) op_1322 (v317[10:0], v163[10:0], v1322[32:0]); // 2.0
    wire [22:0] v1323; shift_adder #(11, 11, 1, 1, 23, 12, 1) op_1323 (v237[10:0], v293[10:0], v1323[22:0]); // 2.0
    wire [12:0] v1324; shift_adder #(11, 12, 1, 1, 13, -1, 1) op_1324 (v234[10:0], v363[11:0], v1324[12:0]); // 2.0
    wire [17:0] v1325; shift_adder #(18, 11, 1, 1, 18, 5, 0) op_1325 (v494[17:0], v386[10:0], v1325[17:0]); // 2.0
    wire [12:0] v1326; shift_adder #(8, 11, 1, 1, 13, 2, 1) op_1326 (v90[7:0], v430[10:0], v1326[12:0]); // 2.0
    wire [12:0] v1327; shift_adder #(12, 12, 1, 1, 13, 1, 0) op_1327 (v495[11:0], v355[11:0], v1327[12:0]); // 2.0
    wire [12:0] v1328; shift_adder #(11, 12, 1, 1, 13, -1, 1) op_1328 (v176[10:0], v304[11:0], v1328[12:0]); // 2.0
    wire [13:0] v1329; shift_adder #(11, 13, 1, 1, 14, -2, 0) op_1329 (v171[10:0], v496[12:0], v1329[13:0]); // 2.0
    wire [14:0] v1330; shift_adder #(11, 14, 1, 1, 15, -4, 0) op_1330 (v212[10:0], v249[13:0], v1330[14:0]); // 2.0
    wire [31:0] v1331; shift_adder #(11, 31, 1, 1, 32, -20, 0) op_1331 (v171[10:0], v381[30:0], v1331[31:0]); // 2.0
    wire [13:0] v1332; shift_adder #(11, 12, 1, 1, 14, -3, 1) op_1332 (v270[10:0], v247[11:0], v1332[13:0]); // 2.0
    wire [11:0] v1333; shift_adder #(11, 11, 1, 1, 12, -1, 0) op_1333 (v133[10:0], v193[10:0], v1333[11:0]); // 2.0
    wire [19:0] v1334; shift_adder #(12, 13, 1, 1, 20, 7, 0) op_1334 (v292[11:0], v272[12:0], v1334[19:0]); // 2.0
    wire [21:0] v1335; shift_adder #(11, 21, 1, 1, 22, -10, 0) op_1335 (v330[10:0], v498[20:0], v1335[21:0]); // 2.0
    wire [12:0] v1336; shift_adder #(8, 11, 1, 1, 13, -4, 0) op_1336 (v101[7:0], v324[10:0], v1336[12:0]); // 2.0
    wire [33:0] v1337; shift_adder #(11, 8, 1, 1, 34, 25, 1) op_1337 (v420[10:0], v126[7:0], v1337[33:0]); // 2.0
    wire [25:0] v1338; shift_adder #(11, 11, 1, 1, 26, 15, 1) op_1338 (v156[10:0], v219[10:0], v1338[25:0]); // 2.0
    wire [13:0] v1339; shift_adder #(14, 12, 1, 1, 14, 1, 0) op_1339 (v499[13:0], v372[11:0], v1339[13:0]); // 2.0
    wire [11:0] v1340; shift_adder #(11, 11, 1, 1, 12, 1, 1) op_1340 (v156[10:0], v177[10:0], v1340[11:0]); // 2.0
    wire [16:0] v1341; shift_adder #(11, 11, 1, 1, 17, 6, 0) op_1341 (v190[10:0], v361[10:0], v1341[16:0]); // 2.0
    wire [21:0] v1342; shift_adder #(11, 11, 1, 1, 22, 11, 0) op_1342 (v193[10:0], v275[10:0], v1342[21:0]); // 2.0
    wire [16:0] v1343; shift_adder #(8, 12, 1, 1, 17, -8, 0) op_1343 (v89[7:0], v500[11:0], v1343[16:0]); // 2.0
    wire [18:0] v1344; shift_adder #(11, 17, 1, 1, 19, -8, 0) op_1344 (v136[10:0], v436[16:0], v1344[18:0]); // 2.0
    wire [21:0] v1345; shift_adder #(19, 10, 1, 1, 22, 12, 0) op_1345 (v376[18:0], v501[9:0], v1345[21:0]); // 2.0
    wire [12:0] v1346; shift_adder #(8, 11, 1, 1, 13, -4, 1) op_1346 (v110[7:0], v141[10:0], v1346[12:0]); // 2.0
    wire [11:0] v1347; shift_adder #(11, 9, 1, 1, 12, -1, 0) op_1347 (v150[10:0], v401[8:0], v1347[11:0]); // 2.0
    wire [11:0] v1348; shift_adder #(12, 9, 1, 1, 12, 1, 0) op_1348 (v502[11:0], v503[8:0], v1348[11:0]); // 2.0
    wire [12:0] v1349; shift_adder #(11, 11, 1, 1, 13, 2, 1) op_1349 (v244[10:0], v289[10:0], v1349[12:0]); // 2.0
    wire [14:0] v1350; shift_adder #(15, 11, 1, 1, 15, 2, 0) op_1350 (v318[14:0], v341[10:0], v1350[14:0]); // 2.0
    wire [14:0] v1351; shift_adder #(11, 11, 1, 1, 15, -4, 0) op_1351 (v136[10:0], v145[10:0], v1351[14:0]); // 2.0
    wire [14:0] v1352; shift_adder #(11, 11, 1, 1, 15, -4, 1) op_1352 (v155[10:0], v135[10:0], v1352[14:0]); // 2.0
    wire [21:0] v1353; shift_adder #(16, 21, 1, 1, 22, -6, 0) op_1353 (v504[15:0], v427[20:0], v1353[21:0]); // 2.0
    wire [29:0] v1354; shift_adder #(11, 11, 1, 1, 30, -19, 0) op_1354 (v175[10:0], v505[10:0], v1354[29:0]); // 2.0
    wire [21:0] v1355; shift_adder #(8, 12, 1, 1, 22, -13, 0) op_1355 (v113[7:0], v164[11:0], v1355[21:0]); // 2.0
    wire [12:0] v1356; shift_adder #(8, 13, 1, 1, 13, -2, 0) op_1356 (v119[7:0], v506[12:0], v1356[12:0]); // 2.0
    wire [13:0] v1357; shift_adder #(13, 11, 1, 1, 14, 2, 0) op_1357 (v416[12:0], v341[10:0], v1357[13:0]); // 2.0
    wire [10:0] v1358; shift_adder #(8, 11, 1, 1, 11, -1, 1) op_1358 (v87[7:0], v195[10:0], v1358[10:0]); // 2.0
    wire [12:0] v1359; shift_adder #(11, 12, 1, 1, 13, 1, 0) op_1359 (v420[10:0], v507[11:0], v1359[12:0]); // 2.0
    wire [15:0] v1360; shift_adder #(8, 12, 1, 1, 16, 4, 0) op_1360 (v87[7:0], v205[11:0], v1360[15:0]); // 2.0
    wire [12:0] v1361; shift_adder #(11, 9, 1, 1, 13, 3, 0) op_1361 (v244[10:0], v508[8:0], v1361[12:0]); // 2.0
    wire [10:0] v1362; shift_adder #(10, 11, 1, 1, 11, 0, 0) op_1362 (v509[9:0], v298[10:0], v1362[10:0]); // 2.0
    wire [10:0] v1363; shift_adder #(10, 10, 1, 1, 11, 0, 0) op_1363 (v466[9:0], v510[9:0], v1363[10:0]); // 2.0
    wire [15:0] v1364; shift_adder #(16, 12, 1, 1, 16, 3, 0) op_1364 (v426[15:0], v224[11:0], v1364[15:0]); // 2.0
    wire [21:0] v1365; shift_adder #(8, 14, 1, 1, 22, 8, 0) op_1365 (v98[7:0], v236[13:0], v1365[21:0]); // 2.0
    wire [36:0] v1366; shift_adder #(35, 9, 1, 1, 37, 27, 0) op_1366 (v511[34:0], v508[8:0], v1366[36:0]); // 2.0
    wire [14:0] v1367; shift_adder #(8, 12, 1, 1, 15, -6, 1) op_1367 (v108[7:0], v304[11:0], v1367[14:0]); // 2.0
    wire [11:0] v1368; shift_adder #(11, 11, 1, 1, 12, 1, 0) op_1368 (v241[10:0], v208[10:0], v1368[11:0]); // 2.0
    wire [29:0] v1369; shift_adder #(8, 11, 1, 1, 30, 19, 0) op_1369 (v95[7:0], v178[10:0], v1369[29:0]); // 2.0
    wire [11:0] v1370; shift_adder #(8, 11, 1, 1, 12, 1, 0) op_1370 (v117[7:0], v294[10:0], v1370[11:0]); // 2.0
    wire [15:0] v1371; shift_adder #(14, 11, 1, 1, 16, 5, 0) op_1371 (v474[13:0], v264[10:0], v1371[15:0]); // 2.0
    wire [11:0] v1372; shift_adder #(11, 11, 1, 1, 12, 0, 1) op_1372 (v132[10:0], v175[10:0], v1372[11:0]); // 2.0
    wire [11:0] v1373; shift_adder #(12, 10, 1, 1, 12, 0, 0) op_1373 (v512[11:0], v466[9:0], v1373[11:0]); // 2.0
    wire [14:0] v1374; shift_adder #(14, 12, 1, 1, 15, 2, 0) op_1374 (v513[13:0], v404[11:0], v1374[14:0]); // 2.0
    wire [12:0] v1375; shift_adder #(8, 11, 1, 1, 13, 2, 1) op_1375 (v81[7:0], v139[10:0], v1375[12:0]); // 2.0
    wire [11:0] v1376; shift_adder #(8, 11, 1, 1, 12, -2, 0) op_1376 (v69[7:0], v275[10:0], v1376[11:0]); // 2.0
    wire [13:0] v1377; shift_adder #(14, 12, 1, 1, 14, 0, 0) op_1377 (v514[13:0], v285[11:0], v1377[13:0]); // 2.0
    wire [13:0] v1378; shift_adder #(11, 11, 1, 1, 14, -3, 1) op_1378 (v283[10:0], v266[10:0], v1378[13:0]); // 2.0
    wire [11:0] v1379; shift_adder #(8, 11, 1, 1, 12, 1, 0) op_1379 (v101[7:0], v210[10:0], v1379[11:0]); // 2.0
    wire [13:0] v1380; shift_adder #(11, 11, 1, 1, 14, 3, 0) op_1380 (v157[10:0], v190[10:0], v1380[13:0]); // 2.0
    wire [13:0] v1381; shift_adder #(8, 11, 1, 1, 14, 3, 0) op_1381 (v115[7:0], v341[10:0], v1381[13:0]); // 2.0
    wire [15:0] v1382; shift_adder #(11, 12, 1, 1, 16, -5, 0) op_1382 (v375[10:0], v183[11:0], v1382[15:0]); // 2.0
    wire [11:0] v1383; shift_adder #(10, 11, 1, 1, 12, -1, 0) op_1383 (v461[9:0], v178[10:0], v1383[11:0]); // 2.0
    wire [19:0] v1384; shift_adder #(8, 12, 1, 1, 20, -11, 1) op_1384 (v118[7:0], v314[11:0], v1384[19:0]); // 2.0
    wire [12:0] v1385; shift_adder #(11, 11, 1, 1, 13, 2, 0) op_1385 (v270[10:0], v341[10:0], v1385[12:0]); // 2.0
    wire [13:0] v1386; shift_adder #(11, 11, 1, 1, 14, -3, 1) op_1386 (v140[10:0], v199[10:0], v1386[13:0]); // 2.0
    wire [14:0] v1387; shift_adder #(11, 11, 1, 1, 15, -4, 1) op_1387 (v323[10:0], v287[10:0], v1387[14:0]); // 2.0
    wire [21:0] v1388; shift_adder #(8, 10, 1, 1, 22, -13, 1) op_1388 (v106[7:0], v516[9:0], v1388[21:0]); // 2.0
    wire [15:0] v1389; shift_adder #(8, 11, 1, 1, 16, 5, 0) op_1389 (v104[7:0], v246[10:0], v1389[15:0]); // 2.0
    wire [25:0] v1390; shift_adder #(10, 26, 1, 1, 26, -12, 0) op_1390 (v428[9:0], v517[25:0], v1390[25:0]); // 2.0
    wire [17:0] v1391; shift_adder #(12, 12, 1, 1, 18, -6, 1) op_1391 (v392[11:0], v392[11:0], v1391[17:0]); // 2.0
    wire [16:0] v1392; shift_adder #(11, 11, 1, 1, 17, 6, 1) op_1392 (v152[10:0], v232[10:0], v1392[16:0]); // 2.0
    wire [12:0] v1393; shift_adder #(11, 11, 1, 1, 13, 2, 1) op_1393 (v234[10:0], v298[10:0], v1393[12:0]); // 2.0
    wire [13:0] v1394; shift_adder #(8, 14, 1, 1, 14, -1, 0) op_1394 (v100[7:0], v499[13:0], v1394[13:0]); // 2.0
    wire [10:0] v1395; shift_adder #(8, 11, 1, 1, 11, -1, 1) op_1395 (v82[7:0], v297[10:0], v1395[10:0]); // 2.0
    wire [24:0] v1396; shift_adder #(10, 10, 1, 1, 25, 15, 1) op_1396 (v510[9:0], v442[9:0], v1396[24:0]); // 2.0
    wire [12:0] v1397; shift_adder #(8, 11, 1, 1, 13, 2, 1) op_1397 (v77[7:0], v136[10:0], v1397[12:0]); // 2.0
    wire [11:0] v1398; shift_adder #(8, 11, 1, 1, 12, -2, 0) op_1398 (v115[7:0], v255[10:0], v1398[11:0]); // 2.0
    wire [11:0] v1399; shift_adder #(11, 11, 1, 1, 12, 1, 1) op_1399 (v276[10:0], v289[10:0], v1399[11:0]); // 2.0
    wire [19:0] v1400; shift_adder #(8, 11, 1, 1, 20, 9, 1) op_1400 (v74[7:0], v215[10:0], v1400[19:0]); // 2.0
    wire [14:0] v1401; shift_adder #(11, 11, 1, 1, 15, 4, 0) op_1401 (v148[10:0], v168[10:0], v1401[14:0]); // 2.0
    wire [15:0] v1402; shift_adder #(14, 9, 1, 1, 16, 6, 0) op_1402 (v472[13:0], v221[8:0], v1402[15:0]); // 2.0
    wire [20:0] v1403; shift_adder #(11, 11, 1, 1, 21, -10, 1) op_1403 (v208[10:0], v518[10:0], v1403[20:0]); // 2.0
    wire [12:0] v1404; shift_adder #(11, 11, 1, 1, 13, -2, 1) op_1404 (v353[10:0], v246[10:0], v1404[12:0]); // 2.0
    wire [24:0] v1405; shift_adder #(11, 11, 1, 1, 25, -14, 1) op_1405 (v250[10:0], v323[10:0], v1405[24:0]); // 2.0
    wire [16:0] v1406; shift_adder #(16, 9, 1, 1, 17, 6, 0) op_1406 (v519[15:0], v369[8:0], v1406[16:0]); // 2.0
    wire [12:0] v1407; shift_adder #(11, 12, 1, 1, 13, -2, 1) op_1407 (v245[10:0], v453[11:0], v1407[12:0]); // 2.0
    wire [11:0] v1408; shift_adder #(11, 11, 1, 1, 12, 1, 0) op_1408 (v317[10:0], v341[10:0], v1408[11:0]); // 2.0
    wire [10:0] v1409; shift_adder #(11, 10, 1, 1, 11, 0, 0) op_1409 (v415[10:0], v520[9:0], v1409[10:0]); // 2.0
    wire [16:0] v1410; shift_adder #(12, 12, 1, 1, 17, -5, 0) op_1410 (v288[11:0], v521[11:0], v1410[16:0]); // 2.0
    wire [19:0] v1411; shift_adder #(11, 12, 1, 1, 20, 8, 1) op_1411 (v297[10:0], v204[11:0], v1411[19:0]); // 2.0
    wire [11:0] v1412; shift_adder #(11, 11, 1, 1, 12, 0, 0) op_1412 (v172[10:0], v455[10:0], v1412[11:0]); // 2.0
    wire [11:0] v1413; shift_adder #(8, 11, 1, 1, 12, -2, 1) op_1413 (v78[7:0], v386[10:0], v1413[11:0]); // 2.0
    wire [15:0] v1414; shift_adder #(11, 11, 1, 1, 16, 5, 1) op_1414 (v188[10:0], v334[10:0], v1414[15:0]); // 2.0
    wire [10:0] v1415; shift_adder #(10, 11, 1, 1, 11, 0, 0) op_1415 (v442[9:0], v163[10:0], v1415[10:0]); // 2.0
    wire [12:0] v1416; shift_adder #(9, 9, 1, 1, 13, -3, 0) op_1416 (v522[8:0], v230[8:0], v1416[12:0]); // 2.0
    wire [14:0] v1417; shift_adder #(11, 11, 1, 1, 15, -4, 0) op_1417 (v218[10:0], v245[10:0], v1417[14:0]); // 2.0
    wire [23:0] v1418; shift_adder #(11, 11, 1, 1, 24, -13, 0) op_1418 (v133[10:0], v299[10:0], v1418[23:0]); // 2.0
    wire [10:0] v1419; shift_adder #(8, 11, 1, 1, 11, -1, 0) op_1419 (v64[7:0], v358[10:0], v1419[10:0]); // 2.0
    wire [13:0] v1420; shift_adder #(8, 11, 1, 1, 14, 3, 0) op_1420 (v69[7:0], v287[10:0], v1420[13:0]); // 2.0
    wire [12:0] v1421; shift_adder #(11, 11, 1, 1, 13, -2, 0) op_1421 (v238[10:0], v268[10:0], v1421[12:0]); // 2.0
    wire [12:0] v1422; shift_adder #(8, 11, 1, 1, 13, -4, 0) op_1422 (v96[7:0], v153[10:0], v1422[12:0]); // 2.0
    wire [18:0] v1423; shift_adder #(11, 12, 1, 1, 19, 7, 0) op_1423 (v172[10:0], v523[11:0], v1423[18:0]); // 2.0
    wire [15:0] v1424; shift_adder #(11, 13, 1, 1, 16, 3, 0) op_1424 (v228[10:0], v524[12:0], v1424[15:0]); // 2.0
    wire [15:0] v1425; shift_adder #(11, 11, 1, 1, 16, 5, 0) op_1425 (v171[10:0], v212[10:0], v1425[15:0]); // 2.0
    wire [10:0] v1426; shift_adder #(8, 11, 1, 1, 11, -1, 0) op_1426 (v110[7:0], v420[10:0], v1426[10:0]); // 2.0
    wire [10:0] v1427; shift_adder #(10, 9, 1, 1, 11, 1, 0) op_1427 (v225[9:0], v479[8:0], v1427[10:0]); // 2.0
    wire [25:0] v1428; shift_adder #(11, 26, 1, 1, 26, -14, 0) op_1428 (v228[10:0], v525[25:0], v1428[25:0]); // 2.0
    wire [14:0] v1429; shift_adder #(8, 12, 1, 1, 15, 3, 1) op_1429 (v102[7:0], v194[11:0], v1429[14:0]); // 2.0
    wire [14:0] v1430; shift_adder #(8, 9, 1, 1, 15, 5, 0) op_1430 (v83[7:0], v370[8:0], v1430[14:0]); // 2.0
    wire [12:0] v1431; shift_adder #(11, 12, 1, 1, 13, -1, 0) op_1431 (v242[10:0], v408[11:0], v1431[12:0]); // 2.0
    wire [32:0] v1432; shift_adder #(10, 8, 1, 1, 33, 24, 1) op_1432 (v446[9:0], v94[7:0], v1432[32:0]); // 2.0
    wire [12:0] v1433; shift_adder #(8, 11, 1, 1, 13, 2, 1) op_1433 (v88[7:0], v276[10:0], v1433[12:0]); // 2.0
    wire [14:0] v1434; shift_adder #(11, 15, 1, 1, 15, -2, 0) op_1434 (v150[10:0], v526[14:0], v1434[14:0]); // 2.0
    wire [36:0] v1435; shift_adder #(10, 11, 1, 1, 37, -27, 1) op_1435 (v459[9:0], v216[10:0], v1435[36:0]); // 2.0
    wire [11:0] v1436; shift_adder #(8, 11, 1, 1, 12, 1, 1) op_1436 (v124[7:0], v320[10:0], v1436[11:0]); // 2.0
    wire [11:0] v1437; shift_adder #(10, 11, 1, 1, 12, -1, 0) op_1437 (v527[9:0], v497[10:0], v1437[11:0]); // 2.0
    wire [12:0] v1438; shift_adder #(8, 11, 1, 1, 13, 2, 0) op_1438 (v102[7:0], v147[10:0], v1438[12:0]); // 2.0
    wire [14:0] v1439; shift_adder #(8, 12, 1, 1, 15, -6, 0) op_1439 (v99[7:0], v174[11:0], v1439[14:0]); // 2.0
    wire [12:0] v1440; shift_adder #(13, 11, 1, 1, 13, 1, 0) op_1440 (v451[12:0], v293[10:0], v1440[12:0]); // 2.0
    wire [32:0] v1441; shift_adder #(12, 15, 1, 1, 33, 18, 0) op_1441 (v292[11:0], v528[14:0], v1441[32:0]); // 2.0
    wire [29:0] v1442; shift_adder #(11, 16, 1, 1, 30, -19, 0) op_1442 (v195[10:0], v166[15:0], v1442[29:0]); // 2.0
    wire [11:0] v1443; shift_adder #(8, 11, 1, 1, 12, -2, 1) op_1443 (v86[7:0], v223[10:0], v1443[11:0]); // 2.0
    wire [24:0] v1444; shift_adder #(11, 11, 1, 1, 25, -14, 1) op_1444 (v155[10:0], v298[10:0], v1444[24:0]); // 2.0
    wire [17:0] v1445; shift_adder #(11, 15, 1, 1, 18, -7, 1) op_1445 (v284[10:0], v253[14:0], v1445[17:0]); // 2.0
    wire [12:0] v1446; shift_adder #(11, 11, 1, 1, 13, -2, 1) op_1446 (v237[10:0], v455[10:0], v1446[12:0]); // 2.0
    wire [15:0] v1447; shift_adder #(11, 11, 1, 1, 16, 5, 0) op_1447 (v172[10:0], v358[10:0], v1447[15:0]); // 2.0
    wire [25:0] v1448; shift_adder #(11, 12, 1, 1, 26, 14, 0) op_1448 (v293[10:0], v214[11:0], v1448[25:0]); // 2.0
    wire [25:0] v1449; shift_adder #(12, 14, 1, 1, 26, 12, 1) op_1449 (v224[11:0], v226[13:0], v1449[25:0]); // 2.0
    wire [23:0] v1450; shift_adder #(24, 11, 1, 1, 24, 10, 0) op_1450 (v529[23:0], v420[10:0], v1450[23:0]); // 2.0
    wire [17:0] v1451; shift_adder #(12, 12, 1, 1, 18, 6, 1) op_1451 (v408[11:0], v521[11:0], v1451[17:0]); // 2.0
    wire [15:0] v1452; shift_adder #(11, 11, 1, 1, 16, -5, 0) op_1452 (v266[10:0], v154[10:0], v1452[15:0]); // 2.0
    wire [17:0] v1453; shift_adder #(11, 11, 1, 1, 18, -7, 0) op_1453 (v157[10:0], v157[10:0], v1453[17:0]); // 2.0
    wire [25:0] v1454; shift_adder #(26, 11, 1, 1, 26, 14, 0) op_1454 (v530[25:0], v270[10:0], v1454[25:0]); // 2.0
    wire [16:0] v1455; shift_adder #(8, 11, 1, 1, 17, -8, 1) op_1455 (v64[7:0], v212[10:0], v1455[16:0]); // 2.0
    wire [12:0] v1456; shift_adder #(11, 11, 1, 1, 13, 2, 1) op_1456 (v328[10:0], v179[10:0], v1456[12:0]); // 2.0
    wire [19:0] v1457; shift_adder #(12, 10, 1, 1, 20, 10, 0) op_1457 (v292[11:0], v468[9:0], v1457[19:0]); // 2.0
    wire [12:0] v1458; shift_adder #(11, 11, 1, 1, 13, -2, 0) op_1458 (v269[10:0], v334[10:0], v1458[12:0]); // 2.0
    wire [12:0] v1459; shift_adder #(11, 11, 1, 1, 13, -2, 0) op_1459 (v297[10:0], v353[10:0], v1459[12:0]); // 2.0
    wire [23:0] v1460; shift_adder #(11, 11, 1, 1, 24, -13, 1) op_1460 (v210[10:0], v153[10:0], v1460[23:0]); // 2.0
    wire [12:0] v1461; shift_adder #(11, 12, 1, 1, 13, 1, 0) op_1461 (v208[10:0], v502[11:0], v1461[12:0]); // 2.0
    wire [11:0] v1462; shift_adder #(11, 11, 1, 1, 12, 0, 0) op_1462 (v200[10:0], v338[10:0], v1462[11:0]); // 2.0
    wire [11:0] v1463; shift_adder #(12, 9, 1, 1, 12, 0, 0) op_1463 (v457[11:0], v309[8:0], v1463[11:0]); // 2.0
    wire [16:0] v1464; shift_adder #(8, 11, 1, 1, 17, -8, 0) op_1464 (v65[7:0], v400[10:0], v1464[16:0]); // 2.0
    wire [10:0] v1465; shift_adder #(11, 9, 1, 1, 11, 0, 0) op_1465 (v203[10:0], v401[8:0], v1465[10:0]); // 2.0
    wire [11:0] v1466; shift_adder #(11, 12, 1, 1, 12, 0, 0) op_1466 (v140[10:0], v453[11:0], v1466[11:0]); // 2.0
    wire [16:0] v1467; shift_adder #(11, 11, 1, 1, 17, 6, 0) op_1467 (v455[10:0], v379[10:0], v1467[16:0]); // 2.0
    wire [11:0] v1468; shift_adder #(11, 11, 1, 1, 12, 1, 1) op_1468 (v203[10:0], v275[10:0], v1468[11:0]); // 2.0
    wire [22:0] v1469; shift_adder #(11, 11, 1, 1, 23, -12, 0) op_1469 (v250[10:0], v140[10:0], v1469[22:0]); // 2.0
    wire [23:0] v1470; shift_adder #(8, 11, 1, 1, 24, -15, 1) op_1470 (v115[7:0], v244[10:0], v1470[23:0]); // 2.0
    wire [12:0] v1471; shift_adder #(11, 12, 1, 1, 13, 1, 0) op_1471 (v181[10:0], v204[11:0], v1471[12:0]); // 2.0
    wire [15:0] v1472; shift_adder #(8, 11, 1, 1, 16, -7, 0) op_1472 (v101[7:0], v218[10:0], v1472[15:0]); // 2.0
    wire [14:0] v1473; shift_adder #(11, 11, 1, 1, 15, 4, 0) op_1473 (v228[10:0], v245[10:0], v1473[14:0]); // 2.0
    wire [22:0] v1474; shift_adder #(11, 12, 1, 1, 23, 11, 1) op_1474 (v156[10:0], v389[11:0], v1474[22:0]); // 2.0
    wire [11:0] v1475; shift_adder #(8, 11, 1, 1, 12, -2, 0) op_1475 (v77[7:0], v362[10:0], v1475[11:0]); // 2.0
    wire [26:0] v1476; shift_adder #(11, 18, 1, 1, 27, -16, 0) op_1476 (v289[10:0], v167[17:0], v1476[26:0]); // 2.0
    wire [14:0] v1477; shift_adder #(8, 11, 1, 1, 15, 4, 1) op_1477 (v126[7:0], v200[10:0], v1477[14:0]); // 2.0
    wire [16:0] v1478; shift_adder #(17, 10, 1, 1, 17, 6, 0) op_1478 (v533[16:0], v510[9:0], v1478[16:0]); // 2.0
    wire [12:0] v1479; shift_adder #(11, 13, 1, 1, 13, -1, 1) op_1479 (v420[10:0], v534[12:0], v1479[12:0]); // 2.0
    wire [13:0] v1480; shift_adder #(11, 13, 1, 1, 14, -3, 0) op_1480 (v443[10:0], v406[12:0], v1480[13:0]); // 2.0
    wire [19:0] v1481; shift_adder #(19, 19, 1, 1, 20, 1, 0) op_1481 (v315[18:0], v536[18:0], v1481[19:0]); // 2.0
    wire [12:0] v1482; shift_adder #(11, 11, 1, 1, 13, 2, 1) op_1482 (v157[10:0], v190[10:0], v1482[12:0]); // 2.0
    wire [25:0] v1483; shift_adder #(8, 11, 1, 1, 26, -17, 0) op_1483 (v74[7:0], v241[10:0], v1483[25:0]); // 2.0
    wire [11:0] v1484; shift_adder #(8, 11, 1, 1, 12, 1, 0) op_1484 (v113[7:0], v269[10:0], v1484[11:0]); // 2.0
    wire [16:0] v1485; shift_adder #(11, 12, 1, 1, 17, 5, 1) op_1485 (v269[10:0], v434[11:0], v1485[16:0]); // 2.0
    wire [25:0] v1486; shift_adder #(25, 9, 1, 1, 26, 16, 0) op_1486 (v537[24:0], v538[8:0], v1486[25:0]); // 2.0
    wire [23:0] v1487; shift_adder #(11, 11, 1, 1, 24, 13, 0) op_1487 (v181[10:0], v172[10:0], v1487[23:0]); // 2.0
    wire [30:0] v1488; shift_adder #(11, 19, 1, 1, 31, -20, 1) op_1488 (v185[10:0], v539[18:0], v1488[30:0]); // 2.0
    wire [35:0] v1489; shift_adder #(12, 9, 1, 1, 36, -24, 1) op_1489 (v159[11:0], v441[8:0], v1489[35:0]); // 2.0
    wire [12:0] v1490; shift_adder #(12, 12, 1, 1, 13, -1, 0) op_1490 (v540[11:0], v541[11:0], v1490[12:0]); // 2.0
    wire [11:0] v1491; shift_adder #(9, 11, 1, 1, 12, -2, 0) op_1491 (v220[8:0], v139[10:0], v1491[11:0]); // 2.0
    wire [10:0] v1492; shift_adder #(8, 11, 1, 1, 11, -1, 0) op_1492 (v66[7:0], v264[10:0], v1492[10:0]); // 2.0
    wire [11:0] v1493; shift_adder #(11, 11, 1, 1, 12, 1, 0) op_1493 (v199[10:0], v345[10:0], v1493[11:0]); // 2.0
    wire [10:0] v1494; shift_adder #(8, 11, 1, 1, 11, -1, 0) op_1494 (v115[7:0], v193[10:0], v1494[10:0]); // 2.0
    wire [12:0] v1495; shift_adder #(10, 11, 1, 1, 13, -2, 0) op_1495 (v542[9:0], v276[10:0], v1495[12:0]); // 2.0
    wire [13:0] v1496; shift_adder #(11, 11, 1, 1, 14, 3, 0) op_1496 (v328[10:0], v238[10:0], v1496[13:0]); // 2.0
    wire [12:0] v1497; shift_adder #(12, 12, 1, 1, 13, 1, 0) op_1497 (v543[11:0], v544[11:0], v1497[12:0]); // 2.0
    wire [11:0] v1498; shift_adder #(11, 11, 1, 1, 12, -1, 1) op_1498 (v188[10:0], v294[10:0], v1498[11:0]); // 2.0
    wire [14:0] v1499; shift_adder #(11, 11, 1, 1, 15, -4, 1) op_1499 (v251[10:0], v293[10:0], v1499[14:0]); // 2.0
    wire [12:0] v1500; shift_adder #(11, 12, 1, 1, 13, -1, 1) op_1500 (v275[10:0], v521[11:0], v1500[12:0]); // 2.0
    wire [12:0] v1501; shift_adder #(13, 11, 1, 1, 13, 0, 0) op_1501 (v272[12:0], v178[10:0], v1501[12:0]); // 2.0
    wire [17:0] v1502; shift_adder #(11, 17, 1, 1, 18, 1, 1) op_1502 (v319[10:0], v545[16:0], v1502[17:0]); // 2.0
    wire [15:0] v1503; shift_adder #(11, 16, 1, 1, 16, -4, 0) op_1503 (v420[10:0], v546[15:0], v1503[15:0]); // 2.0
    wire [27:0] v1504; shift_adder #(12, 11, 1, 1, 28, 17, 1) op_1504 (v243[11:0], v413[10:0], v1504[27:0]); // 2.0
    wire [18:0] v1505; shift_adder #(19, 12, 1, 1, 19, 2, 0) op_1505 (v547[18:0], v151[11:0], v1505[18:0]); // 2.0
    wire [11:0] v1506; shift_adder #(11, 11, 1, 1, 12, 1, 0) op_1506 (v361[10:0], v300[10:0], v1506[11:0]); // 2.0
    wire [13:0] v1507; shift_adder #(12, 10, 1, 1, 14, 4, 1) op_1507 (v383[11:0], v548[9:0], v1507[13:0]); // 2.0
    wire [12:0] v1508; shift_adder #(8, 12, 1, 1, 13, 1, 1) op_1508 (v95[7:0], v333[11:0], v1508[12:0]); // 2.0
    wire [13:0] v1509; shift_adder #(11, 12, 1, 1, 14, 2, 0) op_1509 (v172[10:0], v159[11:0], v1509[13:0]); // 2.0
    wire [17:0] v1510; shift_adder #(11, 11, 1, 1, 18, -7, 1) op_1510 (v284[10:0], v320[10:0], v1510[17:0]); // 2.0
    wire [11:0] v1511; shift_adder #(11, 11, 1, 1, 12, 1, 0) op_1511 (v396[10:0], v393[10:0], v1511[11:0]); // 2.0
    wire [11:0] v1512; shift_adder #(8, 11, 1, 1, 12, -2, 1) op_1512 (v80[7:0], v153[10:0], v1512[11:0]); // 2.0
    wire [13:0] v1513; shift_adder #(8, 11, 1, 1, 14, -5, 0) op_1513 (v126[7:0], v173[10:0], v1513[13:0]); // 2.0
    wire [11:0] v1514; shift_adder #(12, 11, 1, 1, 12, 0, 0) op_1514 (v550[11:0], v242[10:0], v1514[11:0]); // 2.0
    wire [23:0] v1515; shift_adder #(8, 11, 1, 1, 24, -15, 0) op_1515 (v104[7:0], v134[10:0], v1515[23:0]); // 2.0
    wire [13:0] v1516; shift_adder #(11, 11, 1, 1, 14, 3, 0) op_1516 (v145[10:0], v418[10:0], v1516[13:0]); // 2.0
    wire [10:0] v1517; shift_adder #(8, 11, 1, 1, 11, 0, 0) op_1517 (v75[7:0], v287[10:0], v1517[10:0]); // 2.0
    wire [12:0] v1518; shift_adder #(12, 12, 1, 1, 13, 1, 0) op_1518 (v385[11:0], v164[11:0], v1518[12:0]); // 2.0
    wire [16:0] v1519; shift_adder #(11, 17, 1, 1, 17, -5, 1) op_1519 (v259[10:0], v551[16:0], v1519[16:0]); // 2.0
    wire [20:0] v1520; shift_adder #(8, 12, 1, 1, 21, -12, 0) op_1520 (v96[7:0], v325[11:0], v1520[20:0]); // 2.0
    wire [11:0] v1521; shift_adder #(11, 11, 1, 1, 12, 0, 0) op_1521 (v165[10:0], v319[10:0], v1521[11:0]); // 2.0
    wire [13:0] v1522; shift_adder #(11, 12, 1, 1, 14, -3, 1) op_1522 (v241[10:0], v438[11:0], v1522[13:0]); // 2.0
    wire [10:0] v1523; shift_adder #(11, 10, 1, 1, 11, 0, 1) op_1523 (v145[10:0], v450[9:0], v1523[10:0]); // 2.0
    wire [12:0] v1524; shift_adder #(11, 11, 1, 1, 13, 2, 1) op_1524 (v188[10:0], v156[10:0], v1524[12:0]); // 2.0
    wire [15:0] v1525; shift_adder #(11, 11, 1, 1, 16, -5, 0) op_1525 (v294[10:0], v190[10:0], v1525[15:0]); // 2.0
    wire [16:0] v1526; shift_adder #(8, 11, 1, 1, 17, -8, 1) op_1526 (v111[7:0], v178[10:0], v1526[16:0]); // 2.0
    wire [18:0] v1527; shift_adder #(11, 11, 1, 1, 19, 8, 0) op_1527 (v251[10:0], v418[10:0], v1527[18:0]); // 2.0
    wire [27:0] v1528; shift_adder #(8, 11, 1, 1, 28, 17, 1) op_1528 (v108[7:0], v362[10:0], v1528[27:0]); // 2.0
    wire [11:0] v1529; shift_adder #(11, 11, 1, 1, 12, -1, 0) op_1529 (v155[10:0], v152[10:0], v1529[11:0]); // 2.0
    wire [18:0] v1530; shift_adder #(8, 11, 1, 1, 19, -10, 1) op_1530 (v86[7:0], v329[10:0], v1530[18:0]); // 2.0
    wire [15:0] v1531; shift_adder #(11, 11, 1, 1, 16, 5, 0) op_1531 (v297[10:0], v277[10:0], v1531[15:0]); // 2.0
    wire [13:0] v1532; shift_adder #(10, 11, 1, 1, 14, -4, 0) op_1532 (v520[9:0], v233[10:0], v1532[13:0]); // 2.0
    wire [12:0] v1533; shift_adder #(8, 10, 1, 1, 13, -4, 0) op_1533 (v78[7:0], v469[9:0], v1533[12:0]); // 2.0
    wire [11:0] v1534; shift_adder #(8, 11, 1, 1, 12, -2, 0) op_1534 (v91[7:0], v277[10:0], v1534[11:0]); // 2.0
    wire [14:0] v1535; shift_adder #(11, 11, 1, 1, 15, -4, 0) op_1535 (v241[10:0], v396[10:0], v1535[14:0]); // 2.0
    wire [14:0] v1536; shift_adder #(11, 11, 1, 1, 15, -4, 0) op_1536 (v358[10:0], v518[10:0], v1536[14:0]); // 2.0
    wire [11:0] v1537; shift_adder #(8, 11, 1, 1, 12, -3, 1) op_1537 (v112[7:0], v193[10:0], v1537[11:0]); // 2.0
    wire [13:0] v1538; shift_adder #(11, 11, 1, 1, 14, -3, 0) op_1538 (v193[10:0], v217[10:0], v1538[13:0]); // 2.0
    wire [20:0] v1539; shift_adder #(11, 9, 1, 1, 21, 11, 1) op_1539 (v163[10:0], v433[8:0], v1539[20:0]); // 2.0
    wire [16:0] v1540; shift_adder #(11, 11, 1, 1, 17, -6, 1) op_1540 (v270[10:0], v338[10:0], v1540[16:0]); // 2.0
    wire [15:0] v1541; shift_adder #(11, 11, 1, 1, 16, 5, 1) op_1541 (v386[10:0], v367[10:0], v1541[15:0]); // 2.0
    wire [16:0] v1542; shift_adder #(8, 13, 1, 1, 17, -8, 1) op_1542 (v78[7:0], v496[12:0], v1542[16:0]); // 2.0
    wire [10:0] v1543; shift_adder #(10, 9, 1, 1, 11, 1, 0) op_1543 (v554[9:0], v433[8:0], v1543[10:0]); // 2.0
    wire [24:0] v1544; shift_adder #(11, 11, 1, 1, 25, -14, 1) op_1544 (v157[10:0], v393[10:0], v1544[24:0]); // 2.0
    wire [13:0] v1545; shift_adder #(11, 11, 1, 1, 14, -3, 0) op_1545 (v147[10:0], v266[10:0], v1545[13:0]); // 2.0
    wire [16:0] v1546; shift_adder #(11, 11, 1, 1, 17, -6, 1) op_1546 (v148[10:0], v142[10:0], v1546[16:0]); // 2.0
    wire [18:0] v1547; shift_adder #(11, 10, 1, 1, 19, -8, 0) op_1547 (v361[10:0], v428[9:0], v1547[18:0]); // 2.0
    wire [23:0] v1548; shift_adder #(11, 12, 1, 1, 24, 12, 0) op_1548 (v362[10:0], v473[11:0], v1548[23:0]); // 2.0
    wire [13:0] v1549; shift_adder #(11, 14, 1, 1, 14, -2, 0) op_1549 (v300[10:0], v555[13:0], v1549[13:0]); // 2.0
    wire [11:0] v1550; shift_adder #(11, 9, 1, 1, 12, 1, 0) op_1550 (v144[10:0], v556[8:0], v1550[11:0]); // 2.0
    wire [12:0] v1551; shift_adder #(11, 11, 1, 1, 13, 2, 0) op_1551 (v237[10:0], v213[10:0], v1551[12:0]); // 2.0
    wire [15:0] v1552; shift_adder #(8, 11, 1, 1, 16, -7, 0) op_1552 (v111[7:0], v211[10:0], v1552[15:0]); // 2.0
    wire [18:0] v1553; shift_adder #(12, 15, 1, 1, 19, -7, 0) op_1553 (v464[11:0], v557[14:0], v1553[18:0]); // 2.0
    wire [13:0] v1554; shift_adder #(11, 11, 1, 1, 14, -3, 0) op_1554 (v209[10:0], v156[10:0], v1554[13:0]); // 2.0
    wire [11:0] v1555; shift_adder #(11, 11, 1, 1, 12, 1, 0) op_1555 (v218[10:0], v297[10:0], v1555[11:0]); // 2.0
    wire [11:0] v1556; shift_adder #(10, 10, 1, 1, 12, -1, 0) op_1556 (v222[9:0], v450[9:0], v1556[11:0]); // 2.0
    wire [15:0] v1557; shift_adder #(8, 12, 1, 1, 16, 4, 1) op_1557 (v106[7:0], v336[11:0], v1557[15:0]); // 2.0
    wire [11:0] v1558; shift_adder #(8, 10, 1, 1, 12, -3, 1) op_1558 (v124[7:0], v549[9:0], v1558[11:0]); // 2.0
    wire [12:0] v1559; shift_adder #(12, 12, 1, 1, 13, 0, 0) op_1559 (v280[11:0], v447[11:0], v1559[12:0]); // 2.0
    wire [12:0] v1560; shift_adder #(11, 11, 1, 1, 13, -2, 1) op_1560 (v132[10:0], v197[10:0], v1560[12:0]); // 2.0
    wire [17:0] v1561; shift_adder #(11, 12, 1, 1, 18, 6, 1) op_1561 (v324[10:0], v397[11:0], v1561[17:0]); // 2.0
    wire [21:0] v1562; shift_adder #(11, 11, 1, 1, 22, -11, 1) op_1562 (v393[10:0], v329[10:0], v1562[21:0]); // 2.0
    wire [17:0] v1563; shift_adder #(17, 14, 1, 1, 18, 3, 0) op_1563 (v545[16:0], v472[13:0], v1563[17:0]); // 2.0
    wire [15:0] v1564; shift_adder #(11, 11, 1, 1, 16, -5, 0) op_1564 (v245[10:0], v323[10:0], v1564[15:0]); // 2.0
    wire [18:0] v1565; shift_adder #(11, 12, 1, 1, 19, -8, 1) op_1565 (v250[10:0], v372[11:0], v1565[18:0]); // 2.0
    wire [11:0] v1566; shift_adder #(11, 11, 1, 1, 12, -1, 0) op_1566 (v264[10:0], v150[10:0], v1566[11:0]); // 2.0
    wire [19:0] v1567; shift_adder #(8, 11, 1, 1, 20, 9, 0) op_1567 (v93[7:0], v287[10:0], v1567[19:0]); // 2.0
    wire [18:0] v1568; shift_adder #(14, 19, 1, 1, 19, -1, 0) op_1568 (v454[13:0], v558[18:0], v1568[18:0]); // 2.0
    wire [12:0] v1569; shift_adder #(11, 11, 1, 1, 13, -2, 1) op_1569 (v188[10:0], v283[10:0], v1569[12:0]); // 2.0
    wire [11:0] v1570; shift_adder #(11, 11, 1, 1, 12, -1, 1) op_1570 (v162[10:0], v209[10:0], v1570[11:0]); // 2.0
    wire [11:0] v1571; shift_adder #(11, 11, 1, 1, 12, 0, 0) op_1571 (v228[10:0], v223[10:0], v1571[11:0]); // 2.0
    wire [14:0] v1572; shift_adder #(11, 11, 1, 1, 15, -4, 1) op_1572 (v158[10:0], v158[10:0], v1572[14:0]); // 2.0
    wire [11:0] v1573; shift_adder #(8, 11, 1, 1, 12, -2, 1) op_1573 (v120[7:0], v171[10:0], v1573[11:0]); // 2.0
    wire [16:0] v1574; shift_adder #(16, 11, 1, 1, 17, 6, 0) op_1574 (v240[15:0], v266[10:0], v1574[16:0]); // 2.0
    wire [13:0] v1575; shift_adder #(8, 11, 1, 1, 14, 3, 0) op_1575 (v85[7:0], v250[10:0], v1575[13:0]); // 2.0
    wire [14:0] v1576; shift_adder #(11, 11, 1, 1, 15, -4, 0) op_1576 (v264[10:0], v264[10:0], v1576[14:0]); // 2.0
    wire [14:0] v1577; shift_adder #(12, 12, 1, 1, 15, -3, 0) op_1577 (v408[11:0], v305[11:0], v1577[14:0]); // 2.0
    wire [23:0] v1578; shift_adder #(20, 24, 1, 1, 24, -2, 0) op_1578 (v310[19:0], v559[23:0], v1578[23:0]); // 2.0
    wire [26:0] v1579; shift_adder #(11, 13, 1, 1, 27, 14, 0) op_1579 (v229[10:0], v192[12:0], v1579[26:0]); // 2.0
    wire [19:0] v1580; shift_adder #(12, 20, 1, 1, 20, -6, 0) op_1580 (v387[11:0], v560[19:0], v1580[19:0]); // 2.0
    wire [10:0] v1581; shift_adder #(8, 11, 1, 1, 11, -1, 0) op_1581 (v97[7:0], v317[10:0], v1581[10:0]); // 2.0
    wire [12:0] v1582; shift_adder #(12, 11, 1, 1, 13, 1, 0) op_1582 (v512[11:0], v147[10:0], v1582[12:0]); // 2.0
    wire [14:0] v1583; shift_adder #(11, 9, 1, 1, 15, -4, 0) op_1583 (v171[10:0], v490[8:0], v1583[14:0]); // 2.0
    wire [11:0] v1584; shift_adder #(11, 11, 1, 1, 12, 1, 1) op_1584 (v178[10:0], v161[10:0], v1584[11:0]); // 2.0
    wire [11:0] v1585; shift_adder #(11, 11, 1, 1, 12, -1, 1) op_1585 (v136[10:0], v245[10:0], v1585[11:0]); // 2.0
    wire [20:0] v1586; shift_adder #(8, 9, 1, 1, 21, 11, 0) op_1586 (v93[7:0], v561[8:0], v1586[20:0]); // 2.0
    wire [15:0] v1587; shift_adder #(10, 16, 1, 1, 16, -4, 0) op_1587 (v222[9:0], v350[15:0], v1587[15:0]); // 2.0
    wire [12:0] v1588; shift_adder #(11, 11, 1, 1, 13, -2, 0) op_1588 (v375[10:0], v161[10:0], v1588[12:0]); // 2.0
    wire [11:0] v1589; shift_adder #(11, 11, 1, 1, 12, 1, 0) op_1589 (v203[10:0], v216[10:0], v1589[11:0]); // 2.0
    wire [14:0] v1590; shift_adder #(12, 12, 1, 1, 15, 3, 1) op_1590 (v357[11:0], v207[11:0], v1590[14:0]); // 2.0
    wire [12:0] v1591; shift_adder #(11, 10, 1, 1, 13, 3, 0) op_1591 (v255[10:0], v489[9:0], v1591[12:0]); // 2.0
    wire [17:0] v1592; shift_adder #(8, 11, 1, 1, 18, -9, 0) op_1592 (v83[7:0], v142[10:0], v1592[17:0]); // 2.0
    wire [18:0] v1593; shift_adder #(18, 13, 1, 1, 19, 5, 0) op_1593 (v562[17:0], v458[12:0], v1593[18:0]); // 2.0
    wire [12:0] v1594; shift_adder #(12, 11, 1, 1, 13, 1, 0) op_1594 (v321[11:0], v234[10:0], v1594[12:0]); // 2.0
    wire [22:0] v1595; shift_adder #(11, 23, 1, 1, 23, -10, 0) op_1595 (v563[10:0], v564[22:0], v1595[22:0]); // 2.0
    wire [20:0] v1596; shift_adder #(8, 11, 1, 1, 21, -12, 0) op_1596 (v120[7:0], v172[10:0], v1596[20:0]); // 2.0
    wire [33:0] v1597; shift_adder #(8, 11, 1, 1, 34, 23, 1) op_1597 (v83[7:0], v425[10:0], v1597[33:0]); // 2.0
    wire [37:0] v1598; shift_adder #(11, 8, 1, 1, 38, 29, 1) op_1598 (v197[10:0], v88[7:0], v1598[37:0]); // 2.0
    wire [12:0] v1599; shift_adder #(12, 12, 1, 1, 13, -1, 1) op_1599 (v288[11:0], v464[11:0], v1599[12:0]); // 2.0
    wire [11:0] v1600; shift_adder #(11, 11, 1, 1, 12, 1, 0) op_1600 (v210[10:0], v297[10:0], v1600[11:0]); // 2.0
    wire [12:0] v1601; shift_adder #(8, 11, 1, 1, 13, 2, 0) op_1601 (v95[7:0], v237[10:0], v1601[12:0]); // 2.0
    wire [11:0] v1602; shift_adder #(8, 12, 1, 1, 12, -1, 1) op_1602 (v112[7:0], v183[11:0], v1602[11:0]); // 2.0
    wire [19:0] v1603; shift_adder #(8, 18, 1, 1, 20, -11, 1) op_1603 (v72[7:0], v493[17:0], v1603[19:0]); // 2.0
    wire [11:0] v1604; shift_adder #(11, 11, 1, 1, 12, -1, 0) op_1604 (v317[10:0], v299[10:0], v1604[11:0]); // 2.0
    wire [11:0] v1605; shift_adder #(11, 11, 1, 1, 12, 1, 0) op_1605 (v216[10:0], v276[10:0], v1605[11:0]); // 2.0
    wire [15:0] v1606; shift_adder #(11, 16, 1, 1, 16, -4, 0) op_1606 (v324[10:0], v566[15:0], v1606[15:0]); // 2.0
    wire [13:0] v1607; shift_adder #(8, 11, 1, 1, 14, 3, 1) op_1607 (v121[7:0], v232[10:0], v1607[13:0]); // 2.0
    wire [12:0] v1608; shift_adder #(10, 11, 1, 1, 13, -3, 0) op_1608 (v567[9:0], v175[10:0], v1608[12:0]); // 2.0
    wire [14:0] v1609; shift_adder #(11, 14, 1, 1, 15, 1, 1) op_1609 (v238[10:0], v342[13:0], v1609[14:0]); // 2.0
    wire [13:0] v1610; shift_adder #(11, 12, 1, 1, 14, 2, 1) op_1610 (v284[10:0], v184[11:0], v1610[13:0]); // 2.0
    wire [14:0] v1611; shift_adder #(11, 11, 1, 1, 15, 4, 1) op_1611 (v216[10:0], v374[10:0], v1611[14:0]); // 2.0
    wire [11:0] v1612; shift_adder #(8, 9, 1, 1, 12, 2, 0) op_1612 (v64[7:0], v561[8:0], v1612[11:0]); // 2.0
    wire [10:0] v1613; shift_adder #(11, 9, 1, 1, 11, 0, 0) op_1613 (v200[10:0], v568[8:0], v1613[10:0]); // 2.0
    wire [11:0] v1614; shift_adder #(9, 11, 1, 1, 12, -2, 0) op_1614 (v405[8:0], v281[10:0], v1614[11:0]); // 2.0
    wire [10:0] v1615; shift_adder #(10, 11, 1, 1, 11, 0, 0) op_1615 (v569[9:0], v208[10:0], v1615[10:0]); // 2.0
    wire [12:0] v1616; shift_adder #(11, 11, 1, 1, 13, 2, 0) op_1616 (v139[10:0], v338[10:0], v1616[12:0]); // 2.0
    wire [16:0] v1617; shift_adder #(11, 17, 1, 1, 17, -5, 0) op_1617 (v152[10:0], v143[16:0], v1617[16:0]); // 2.0
    wire [16:0] v1618; shift_adder #(8, 11, 1, 1, 17, -8, 0) op_1618 (v68[7:0], v208[10:0], v1618[16:0]); // 2.0
    wire [16:0] v1619; shift_adder #(8, 11, 1, 1, 17, 6, 1) op_1619 (v104[7:0], v195[10:0], v1619[16:0]); // 2.0
    wire [15:0] v1620; shift_adder #(11, 11, 1, 1, 16, 5, 0) op_1620 (v238[10:0], v172[10:0], v1620[15:0]); // 2.0
    wire [12:0] v1621; shift_adder #(8, 12, 1, 1, 13, -3, 1) op_1621 (v99[7:0], v325[11:0], v1621[12:0]); // 2.0
    wire [23:0] v1622; shift_adder #(11, 11, 1, 1, 24, 13, 0) op_1622 (v136[10:0], v289[10:0], v1622[23:0]); // 2.0
    wire [13:0] v1623; shift_adder #(11, 13, 1, 1, 14, -3, 0) op_1623 (v208[10:0], v496[12:0], v1623[13:0]); // 2.0
    wire [16:0] v1624; shift_adder #(11, 17, 1, 1, 17, -4, 0) op_1624 (v570[10:0], v533[16:0], v1624[16:0]); // 2.0
    wire [24:0] v1625; shift_adder #(8, 10, 1, 1, 25, -16, 0) op_1625 (v83[7:0], v225[9:0], v1625[24:0]); // 2.0
    wire [18:0] v1626; shift_adder #(11, 11, 1, 1, 19, 8, 1) op_1626 (v156[10:0], v420[10:0], v1626[18:0]); // 2.0
    wire [10:0] v1627; shift_adder #(8, 10, 1, 1, 11, -2, 1) op_1627 (v110[7:0], v170[9:0], v1627[10:0]); // 2.0
    wire [14:0] v1628; shift_adder #(11, 12, 1, 1, 15, 3, 1) op_1628 (v223[10:0], v137[11:0], v1628[14:0]); // 2.0
    wire [14:0] v1629; shift_adder #(11, 11, 1, 1, 15, 4, 1) op_1629 (v277[10:0], v246[10:0], v1629[14:0]); // 2.0
    wire [15:0] v1630; shift_adder #(13, 14, 1, 1, 16, 2, 0) op_1630 (v344[12:0], v571[13:0], v1630[15:0]); // 2.0
    wire [11:0] v1631; shift_adder #(11, 12, 1, 1, 12, 0, 0) op_1631 (v374[10:0], v183[11:0], v1631[11:0]); // 2.0
    wire [14:0] v1632; shift_adder #(12, 12, 1, 1, 15, -3, 0) op_1632 (v227[11:0], v333[11:0], v1632[14:0]); // 2.0
    wire [12:0] v1633; shift_adder #(10, 9, 1, 1, 13, 3, 0) op_1633 (v572[9:0], v401[8:0], v1633[12:0]); // 2.0
    wire [24:0] v1634; shift_adder #(11, 11, 1, 1, 25, -14, 0) op_1634 (v338[10:0], v213[10:0], v1634[24:0]); // 2.0
    wire [21:0] v1635; shift_adder #(11, 13, 1, 1, 22, -11, 0) op_1635 (v244[10:0], v416[12:0], v1635[21:0]); // 2.0
    wire [10:0] v1636; shift_adder #(8, 11, 1, 1, 11, 0, 1) op_1636 (v89[7:0], v199[10:0], v1636[10:0]); // 2.0
    wire [11:0] v1637; shift_adder #(11, 11, 1, 1, 12, -1, 0) op_1637 (v210[10:0], v367[10:0], v1637[11:0]); // 2.0
    wire [10:0] v1638; shift_adder #(11, 9, 1, 1, 11, 0, 0) op_1638 (v215[10:0], v531[8:0], v1638[10:0]); // 2.0
    wire [12:0] v1639; shift_adder #(9, 11, 1, 1, 13, 2, 0) op_1639 (v395[8:0], v283[10:0], v1639[12:0]); // 2.0
    wire [11:0] v1640; shift_adder #(11, 9, 1, 1, 12, 1, 0) op_1640 (v574[10:0], v575[8:0], v1640[11:0]); // 2.0
    wire [11:0] v1641; shift_adder #(11, 10, 1, 1, 12, 1, 0) op_1641 (v162[10:0], v445[9:0], v1641[11:0]); // 2.0
    wire [11:0] v1642; shift_adder #(11, 11, 1, 1, 12, -1, 1) op_1642 (v320[10:0], v259[10:0], v1642[11:0]); // 2.0
    wire [18:0] v1643; shift_adder #(11, 11, 1, 1, 19, 8, 1) op_1643 (v162[10:0], v142[10:0], v1643[18:0]); // 2.0
    wire [18:0] v1644; shift_adder #(11, 11, 1, 1, 19, -8, 0) op_1644 (v152[10:0], v293[10:0], v1644[18:0]); // 2.0
    wire [22:0] v1645; shift_adder #(11, 11, 1, 1, 23, -12, 0) op_1645 (v334[10:0], v358[10:0], v1645[22:0]); // 2.0
    wire [36:0] v1646; shift_adder #(12, 8, 1, 1, 37, 28, 1) op_1646 (v292[11:0], v81[7:0], v1646[36:0]); // 2.0
    wire [11:0] v1647; shift_adder #(10, 11, 1, 1, 12, -1, 0) op_1647 (v576[9:0], v134[10:0], v1647[11:0]); // 2.0
    wire [22:0] v1648; shift_adder #(8, 11, 1, 1, 23, -14, 0) op_1648 (v127[7:0], v232[10:0], v1648[22:0]); // 2.0
    wire [11:0] v1649; shift_adder #(10, 11, 1, 1, 12, 1, 0) op_1649 (v548[9:0], v577[10:0], v1649[11:0]); // 2.0
    wire [17:0] v1650; shift_adder #(8, 11, 1, 1, 18, -9, 0) op_1650 (v124[7:0], v375[10:0], v1650[17:0]); // 2.0
    wire [11:0] v1651; shift_adder #(11, 10, 1, 1, 12, 1, 0) op_1651 (v181[10:0], v569[9:0], v1651[11:0]); // 2.0
    wire [19:0] v1652; shift_adder #(11, 11, 1, 1, 20, 9, 0) op_1652 (v251[10:0], v219[10:0], v1652[19:0]); // 2.0
    wire [28:0] v1653; shift_adder #(11, 11, 1, 1, 29, 18, 1) op_1653 (v319[10:0], v169[10:0], v1653[28:0]); // 2.0
    wire [31:0] v1654; shift_adder #(8, 9, 1, 1, 32, 22, 0) op_1654 (v81[7:0], v490[8:0], v1654[31:0]); // 2.0
    wire [11:0] v1655; shift_adder #(11, 9, 1, 1, 12, 2, 0) op_1655 (v255[10:0], v322[8:0], v1655[11:0]); // 2.0
    wire [21:0] v1656; shift_adder #(20, 13, 1, 1, 22, 9, 0) op_1656 (v484[19:0], v578[12:0], v1656[21:0]); // 2.0
    wire [26:0] v1657; shift_adder #(8, 11, 1, 1, 27, 16, 0) op_1657 (v66[7:0], v136[10:0], v1657[26:0]); // 2.0
    wire [11:0] v1658; shift_adder #(11, 10, 1, 1, 12, -1, 0) op_1658 (v210[10:0], v446[9:0], v1658[11:0]); // 2.0
    wire [11:0] v1659; shift_adder #(11, 11, 1, 1, 12, 0, 1) op_1659 (v190[10:0], v297[10:0], v1659[11:0]); // 2.0
    wire [12:0] v1660; shift_adder #(8, 11, 1, 1, 13, 2, 0) op_1660 (v117[7:0], v430[10:0], v1660[12:0]); // 2.0
    wire [12:0] v1661; shift_adder #(11, 11, 1, 1, 13, 2, 1) op_1661 (v156[10:0], v234[10:0], v1661[12:0]); // 2.0
    wire [22:0] v1662; shift_adder #(11, 14, 1, 1, 23, 9, 0) op_1662 (v175[10:0], v488[13:0], v1662[22:0]); // 2.0
    wire [26:0] v1663; shift_adder #(12, 25, 1, 1, 27, -15, 0) op_1663 (v579[11:0], v261[24:0], v1663[26:0]); // 2.0
    wire [21:0] v1664; shift_adder #(11, 9, 1, 1, 22, -11, 1) op_1664 (v287[10:0], v316[8:0], v1664[21:0]); // 2.0
    wire [12:0] v1665; shift_adder #(11, 11, 1, 1, 13, 2, 0) op_1665 (v215[10:0], v418[10:0], v1665[12:0]); // 2.0
    wire [19:0] v1666; shift_adder #(11, 15, 1, 1, 20, 5, 1) op_1666 (v212[10:0], v313[14:0], v1666[19:0]); // 2.0
    wire [24:0] v1667; shift_adder #(11, 11, 1, 1, 25, 14, 1) op_1667 (v246[10:0], v352[10:0], v1667[24:0]); // 2.0
    wire [22:0] v1668; shift_adder #(23, 11, 1, 1, 23, 5, 0) op_1668 (v580[22:0], v581[10:0], v1668[22:0]); // 2.0
    wire [11:0] v1669; shift_adder #(8, 11, 1, 1, 12, -3, 1) op_1669 (v111[7:0], v153[10:0], v1669[11:0]); // 2.0
    wire [12:0] v1670; shift_adder #(11, 11, 1, 1, 13, -2, 0) op_1670 (v158[10:0], v264[10:0], v1670[12:0]); // 2.0
    wire [21:0] v1671; shift_adder #(8, 9, 1, 1, 22, 12, 0) op_1671 (v114[7:0], v395[8:0], v1671[21:0]); // 2.0
    wire [15:0] v1672; shift_adder #(12, 15, 1, 1, 16, -3, 0) op_1672 (v582[11:0], v295[14:0], v1672[15:0]); // 2.0
    wire [13:0] v1673; shift_adder #(11, 14, 1, 1, 14, -2, 0) op_1673 (v153[10:0], v417[13:0], v1673[13:0]); // 2.0
    wire [16:0] v1674; shift_adder #(11, 11, 1, 1, 17, 6, 0) op_1674 (v251[10:0], v242[10:0], v1674[16:0]); // 2.0
    wire [17:0] v1675; shift_adder #(9, 16, 1, 1, 18, -8, 0) op_1675 (v401[8:0], v583[15:0], v1675[17:0]); // 2.0
    wire [13:0] v1676; shift_adder #(11, 11, 1, 1, 14, -3, 0) op_1676 (v518[10:0], v150[10:0], v1676[13:0]); // 2.0
    wire [12:0] v1677; shift_adder #(12, 12, 1, 1, 13, 1, 0) op_1677 (v365[11:0], v398[11:0], v1677[12:0]); // 2.0
    wire [13:0] v1678; shift_adder #(11, 11, 1, 1, 14, 3, 0) op_1678 (v233[10:0], v187[10:0], v1678[13:0]); // 2.0
    wire [13:0] v1679; shift_adder #(11, 11, 1, 1, 14, 3, 0) op_1679 (v293[10:0], v213[10:0], v1679[13:0]); // 2.0
    wire [13:0] v1680; shift_adder #(11, 14, 1, 1, 14, -1, 0) op_1680 (v241[10:0], v394[13:0], v1680[13:0]); // 2.0
    wire [14:0] v1681; shift_adder #(8, 11, 1, 1, 15, -6, 1) op_1681 (v92[7:0], v178[10:0], v1681[14:0]); // 2.0
    wire [15:0] v1682; shift_adder #(8, 11, 1, 1, 16, 5, 1) op_1682 (v103[7:0], v268[10:0], v1682[15:0]); // 2.0
    wire [19:0] v1683; shift_adder #(16, 10, 1, 1, 20, 10, 0) op_1683 (v390[15:0], v584[9:0], v1683[19:0]); // 2.0
    wire [16:0] v1684; shift_adder #(14, 15, 1, 1, 17, -3, 1) op_1684 (v236[13:0], v253[14:0], v1684[16:0]); // 2.0
    wire [22:0] v1685; shift_adder #(11, 10, 1, 1, 23, 13, 1) op_1685 (v209[10:0], v459[9:0], v1685[22:0]); // 2.0
    wire [11:0] v1686; shift_adder #(11, 11, 1, 1, 12, 1, 1) op_1686 (v245[10:0], v303[10:0], v1686[11:0]); // 2.0
    wire [26:0] v1687; shift_adder #(11, 11, 1, 1, 27, -16, 0) op_1687 (v269[10:0], v343[10:0], v1687[26:0]); // 2.0
    wire [14:0] v1688; shift_adder #(11, 12, 1, 1, 15, -4, 0) op_1688 (v175[10:0], v392[11:0], v1688[14:0]); // 2.0
    wire [11:0] v1689; shift_adder #(11, 11, 1, 1, 12, 1, 0) op_1689 (v298[10:0], v386[10:0], v1689[11:0]); // 2.0
    wire [14:0] v1690; shift_adder #(12, 12, 1, 1, 15, 3, 1) op_1690 (v333[11:0], v304[11:0], v1690[14:0]); // 2.0
    wire [15:0] v1691; shift_adder #(12, 10, 1, 1, 16, 6, 0) op_1691 (v337[11:0], v585[9:0], v1691[15:0]); // 2.0
    wire [17:0] v1692; shift_adder #(11, 11, 1, 1, 18, -7, 0) op_1692 (v141[10:0], v199[10:0], v1692[17:0]); // 2.0
    wire [30:0] v1693; shift_adder #(11, 14, 1, 1, 31, 17, 1) op_1693 (v216[10:0], v249[13:0], v1693[30:0]); // 2.0
    wire [11:0] v1694; shift_adder #(8, 11, 1, 1, 12, 1, 0) op_1694 (v100[7:0], v212[10:0], v1694[11:0]); // 2.0
    wire [13:0] v1695; shift_adder #(11, 11, 1, 1, 14, 3, 1) op_1695 (v386[10:0], v133[10:0], v1695[13:0]); // 2.0
    wire [12:0] v1696; shift_adder #(11, 11, 1, 1, 13, -2, 1) op_1696 (v238[10:0], v206[10:0], v1696[12:0]); // 2.0
    wire [19:0] v1697; shift_adder #(12, 11, 1, 1, 20, 9, 0) op_1697 (v333[11:0], v374[10:0], v1697[19:0]); // 2.0
    wire [27:0] v1698; shift_adder #(12, 12, 1, 1, 28, -16, 0) op_1698 (v288[11:0], v586[11:0], v1698[27:0]); // 2.0
    wire [27:0] v1699; shift_adder #(19, 22, 1, 1, 28, -9, 1) op_1699 (v376[18:0], v587[21:0], v1699[27:0]); // 2.0
    wire [16:0] v1700; shift_adder #(11, 11, 1, 1, 17, -6, 0) op_1700 (v152[10:0], v217[10:0], v1700[16:0]); // 2.0
    wire [18:0] v1701; shift_adder #(9, 10, 1, 1, 19, 9, 0) op_1701 (v316[8:0], v527[9:0], v1701[18:0]); // 2.0
    wire [33:0] v1702; shift_adder #(12, 34, 1, 1, 34, -21, 0) op_1702 (v475[11:0], v588[33:0], v1702[33:0]); // 2.0
    wire [23:0] v1703; shift_adder #(15, 12, 1, 1, 24, -9, 1) op_1703 (v253[14:0], v385[11:0], v1703[23:0]); // 2.0
    wire [12:0] v1704; shift_adder #(8, 11, 1, 1, 13, 2, 1) op_1704 (v122[7:0], v211[10:0], v1704[12:0]); // 2.0
    wire [13:0] v1705; shift_adder #(12, 10, 1, 1, 14, 4, 0) op_1705 (v589[11:0], v549[9:0], v1705[13:0]); // 2.0
    wire [12:0] v1706; shift_adder #(12, 12, 1, 1, 13, 0, 0) op_1706 (v544[11:0], v194[11:0], v1706[12:0]); // 2.0
    wire [32:0] v1707; shift_adder #(14, 32, 1, 1, 33, -18, 0) op_1707 (v590[13:0], v591[31:0], v1707[32:0]); // 2.0
    wire [11:0] v1708; shift_adder #(11, 12, 1, 1, 12, 0, 1) op_1708 (v132[10:0], v137[11:0], v1708[11:0]); // 2.0
    wire [17:0] v1709; shift_adder #(9, 13, 1, 1, 18, -8, 0) op_1709 (v322[8:0], v296[12:0], v1709[17:0]); // 2.0
    wire [27:0] v1710; shift_adder #(11, 15, 1, 1, 28, -17, 1) op_1710 (v158[10:0], v471[14:0], v1710[27:0]); // 2.0
    wire [10:0] v1711; shift_adder #(8, 11, 1, 1, 11, -1, 0) op_1711 (v79[7:0], v242[10:0], v1711[10:0]); // 2.0
    wire [27:0] v1712; shift_adder #(9, 28, 1, 1, 28, -18, 0) op_1712 (v368[8:0], v593[27:0], v1712[27:0]); // 2.0
    wire [11:0] v1713; shift_adder #(11, 9, 1, 1, 12, 1, 0) op_1713 (v206[10:0], v370[8:0], v1713[11:0]); // 2.0
    wire [20:0] v1714; shift_adder #(11, 11, 1, 1, 21, 10, 0) op_1714 (v133[10:0], v303[10:0], v1714[20:0]); // 2.0
    wire [17:0] v1715; shift_adder #(8, 11, 1, 1, 18, 7, 1) op_1715 (v76[7:0], v264[10:0], v1715[17:0]); // 2.0
    wire [16:0] v1716; shift_adder #(16, 9, 1, 1, 17, 6, 1) op_1716 (v426[15:0], v369[8:0], v1716[16:0]); // 2.0
    wire [15:0] v1717; shift_adder #(11, 11, 1, 1, 16, -5, 0) op_1717 (v251[10:0], v298[10:0], v1717[15:0]); // 2.0
    wire [13:0] v1718; shift_adder #(11, 11, 1, 1, 14, -3, 0) op_1718 (v153[10:0], v301[10:0], v1718[13:0]); // 2.0
    wire [15:0] v1719; shift_adder #(11, 11, 1, 1, 16, -5, 0) op_1719 (v211[10:0], v201[10:0], v1719[15:0]); // 2.0
    wire [12:0] v1720; shift_adder #(11, 12, 1, 1, 13, -2, 0) op_1720 (v237[10:0], v579[11:0], v1720[12:0]); // 2.0
    wire [14:0] v1721; shift_adder #(11, 14, 1, 1, 15, 1, 1) op_1721 (v455[10:0], v236[13:0], v1721[14:0]); // 2.0
    wire [20:0] v1722; shift_adder #(8, 15, 1, 1, 21, -12, 0) op_1722 (v78[7:0], v431[14:0], v1722[20:0]); // 2.0
    wire [14:0] v1723; shift_adder #(12, 10, 1, 1, 15, 5, 0) op_1723 (v184[11:0], v446[9:0], v1723[14:0]); // 2.0
    wire [13:0] v1724; shift_adder #(11, 11, 1, 1, 14, -3, 0) op_1724 (v250[10:0], v276[10:0], v1724[13:0]); // 2.0
    wire [11:0] v1725; shift_adder #(11, 11, 1, 1, 12, -1, 0) op_1725 (v375[10:0], v218[10:0], v1725[11:0]); // 2.0
    wire [11:0] v1726; shift_adder #(11, 11, 1, 1, 12, 1, 1) op_1726 (v173[10:0], v208[10:0], v1726[11:0]); // 2.0
    wire [28:0] v1727; shift_adder #(8, 16, 1, 1, 29, 13, 1) op_1727 (v67[7:0], v594[15:0], v1727[28:0]); // 2.0
    wire [14:0] v1728; shift_adder #(12, 14, 1, 1, 15, -3, 0) op_1728 (v423[11:0], v460[13:0], v1728[14:0]); // 2.0
    wire [23:0] v1729; shift_adder #(8, 10, 1, 1, 24, 14, 1) op_1729 (v123[7:0], v461[9:0], v1729[23:0]); // 2.0
    wire [11:0] v1730; shift_adder #(8, 11, 1, 1, 12, -3, 0) op_1730 (v73[7:0], v161[10:0], v1730[11:0]); // 2.0
    wire [24:0] v1731; shift_adder #(11, 25, 1, 1, 25, -13, 0) op_1731 (v238[10:0], v595[24:0], v1731[24:0]); // 2.0
    wire [24:0] v1732; shift_adder #(11, 12, 1, 1, 25, -14, 0) op_1732 (v171[10:0], v372[11:0], v1732[24:0]); // 2.0
    wire [22:0] v1733; shift_adder #(11, 11, 1, 1, 23, -12, 0) op_1733 (v251[10:0], v264[10:0], v1733[22:0]); // 2.0
    wire [23:0] v1734; shift_adder #(8, 11, 1, 1, 24, 13, 0) op_1734 (v120[7:0], v299[10:0], v1734[23:0]); // 2.0
    wire [16:0] v1735; shift_adder #(10, 16, 1, 1, 17, -7, 0) op_1735 (v509[9:0], v596[15:0], v1735[16:0]); // 2.0
    wire [12:0] v1736; shift_adder #(11, 11, 1, 1, 13, 2, 1) op_1736 (v144[10:0], v142[10:0], v1736[12:0]); // 2.0
    wire [13:0] v1737; shift_adder #(12, 11, 1, 1, 14, -2, 0) op_1737 (v521[11:0], v218[10:0], v1737[13:0]); // 2.0
    wire [14:0] v1738; shift_adder #(11, 11, 1, 1, 15, 4, 1) op_1738 (v269[10:0], v358[10:0], v1738[14:0]); // 2.0
    wire [19:0] v1739; shift_adder #(17, 12, 1, 1, 20, 8, 0) op_1739 (v436[16:0], v288[11:0], v1739[19:0]); // 2.0
    wire [14:0] v1740; shift_adder #(11, 13, 1, 1, 15, 2, 0) op_1740 (v301[10:0], v192[12:0], v1740[14:0]); // 2.0
    wire [12:0] v1741; shift_adder #(11, 12, 1, 1, 13, -2, 1) op_1741 (v352[10:0], v408[11:0], v1741[12:0]); // 2.0
    wire [10:0] v1742; shift_adder #(9, 11, 1, 1, 11, 0, 0) op_1742 (v368[8:0], v215[10:0], v1742[10:0]); // 2.0
    wire [22:0] v1743; shift_adder #(11, 9, 1, 1, 23, 14, 1) op_1743 (v268[10:0], v360[8:0], v1743[22:0]); // 2.0
    wire [23:0] v1744; shift_adder #(22, 16, 1, 1, 24, 8, 0) op_1744 (v587[21:0], v166[15:0], v1744[23:0]); // 2.0
    wire [11:0] v1745; shift_adder #(11, 11, 1, 1, 12, -1, 1) op_1745 (v190[10:0], v209[10:0], v1745[11:0]); // 2.0
    wire [29:0] v1746; shift_adder #(11, 12, 1, 1, 30, 18, 0) op_1746 (v375[10:0], v372[11:0], v1746[29:0]); // 2.0
    wire [20:0] v1747; shift_adder #(11, 19, 1, 1, 21, -10, 0) op_1747 (v301[10:0], v597[18:0], v1747[20:0]); // 2.0
    wire [18:0] v1748; shift_adder #(8, 12, 1, 1, 19, 7, 0) op_1748 (v69[7:0], v204[11:0], v1748[18:0]); // 2.0
    wire [13:0] v1749; shift_adder #(11, 11, 1, 1, 14, -3, 1) op_1749 (v181[10:0], v193[10:0], v1749[13:0]); // 2.0
    wire [17:0] v1750; shift_adder #(9, 13, 1, 1, 18, -8, 0) op_1750 (v128[8:0], v598[12:0], v1750[17:0]); // 2.0
    wire [25:0] v1751; shift_adder #(11, 21, 1, 1, 26, -15, 1) op_1751 (v157[10:0], v599[20:0], v1751[25:0]); // 2.0
    wire [11:0] v1752; shift_adder #(11, 11, 1, 1, 12, 1, 1) op_1752 (v518[10:0], v600[10:0], v1752[11:0]); // 2.0
    wire [23:0] v1753; shift_adder #(11, 11, 1, 1, 24, 13, 0) op_1753 (v219[10:0], v300[10:0], v1753[23:0]); // 2.0
    wire [11:0] v1754; shift_adder #(8, 11, 1, 1, 12, -2, 1) op_1754 (v77[7:0], v341[10:0], v1754[11:0]); // 2.0
    wire [21:0] v1755; shift_adder #(9, 20, 1, 1, 22, -12, 0) op_1755 (v531[8:0], v484[19:0], v1755[21:0]); // 2.0
    wire [11:0] v1756; shift_adder #(11, 11, 1, 1, 12, 0, 1) op_1756 (v229[10:0], v352[10:0], v1756[11:0]); // 2.0
    wire [11:0] v1757; shift_adder #(10, 11, 1, 1, 12, -1, 0) op_1757 (v469[9:0], v213[10:0], v1757[11:0]); // 2.0
    wire [11:0] v1758; shift_adder #(11, 12, 1, 1, 12, 0, 0) op_1758 (v199[10:0], v383[11:0], v1758[11:0]); // 2.0
    wire [12:0] v1759; shift_adder #(13, 11, 1, 1, 13, 1, 0) op_1759 (v601[12:0], v173[10:0], v1759[12:0]); // 2.0
    wire [21:0] v1760; shift_adder #(12, 11, 1, 1, 22, 11, 0) op_1760 (v336[11:0], v281[10:0], v1760[21:0]); // 2.0
    wire [11:0] v1761; shift_adder #(11, 11, 1, 1, 12, -1, 0) op_1761 (v487[10:0], v602[10:0], v1761[11:0]); // 2.0
    wire [15:0] v1762; shift_adder #(11, 11, 1, 1, 16, 5, 0) op_1762 (v206[10:0], v284[10:0], v1762[15:0]); // 2.0
    wire [29:0] v1763; shift_adder #(20, 30, 1, 1, 30, -5, 0) op_1763 (v604[19:0], v605[29:0], v1763[29:0]); // 2.0
    wire [18:0] v1764; shift_adder #(8, 11, 1, 1, 19, 8, 0) op_1764 (v66[7:0], v251[10:0], v1764[18:0]); // 2.0
    wire [11:0] v1765; shift_adder #(10, 11, 1, 1, 12, 1, 0) op_1765 (v606[9:0], v242[10:0], v1765[11:0]); // 2.0
    wire [12:0] v1766; shift_adder #(11, 11, 1, 1, 13, 2, 0) op_1766 (v607[10:0], v208[10:0], v1766[12:0]); // 2.0
    wire [14:0] v1767; shift_adder #(11, 11, 1, 1, 15, -4, 1) op_1767 (v301[10:0], v396[10:0], v1767[14:0]); // 2.0
    wire [33:0] v1768; shift_adder #(33, 10, 1, 1, 34, 23, 0) op_1768 (v608[32:0], v609[9:0], v1768[33:0]); // 2.0
    wire [14:0] v1769; shift_adder #(8, 10, 1, 1, 15, 5, 0) op_1769 (v79[7:0], v610[9:0], v1769[14:0]); // 2.0
    wire [24:0] v1770; shift_adder #(11, 25, 1, 1, 25, -10, 0) op_1770 (v396[10:0], v611[24:0], v1770[24:0]); // 2.0
    wire [27:0] v1771; shift_adder #(8, 11, 1, 1, 28, 17, 1) op_1771 (v78[7:0], v329[10:0], v1771[27:0]); // 2.0
    wire [18:0] v1772; shift_adder #(11, 13, 1, 1, 19, -8, 0) op_1772 (v245[10:0], v346[12:0], v1772[18:0]); // 2.0
    wire [32:0] v1773; shift_adder #(8, 25, 1, 1, 33, -24, 0) op_1773 (v65[7:0], v595[24:0], v1773[32:0]); // 2.0
    wire [14:0] v1774; shift_adder #(11, 11, 1, 1, 15, 4, 0) op_1774 (v210[10:0], v455[10:0], v1774[14:0]); // 2.0
    wire [11:0] v1775; shift_adder #(11, 11, 1, 1, 12, 1, 0) op_1775 (v300[10:0], v612[10:0], v1775[11:0]); // 2.0
    wire [11:0] v1776; shift_adder #(9, 12, 1, 1, 12, 0, 0) op_1776 (v220[8:0], v462[11:0], v1776[11:0]); // 2.0
    wire [27:0] v1777; shift_adder #(27, 12, 1, 1, 28, 16, 0) op_1777 (v613[26:0], v614[11:0], v1777[27:0]); // 2.0
    wire [17:0] v1778; shift_adder #(11, 17, 1, 1, 18, 1, 1) op_1778 (v155[10:0], v615[16:0], v1778[17:0]); // 2.0
    wire [32:0] v1779; shift_adder #(12, 14, 1, 1, 33, -21, 0) op_1779 (v423[11:0], v483[13:0], v1779[32:0]); // 2.0
    wire [14:0] v1780; shift_adder #(10, 15, 1, 1, 15, -4, 0) op_1780 (v291[9:0], v456[14:0], v1780[14:0]); // 2.0
    wire [12:0] v1781; shift_adder #(11, 12, 1, 1, 13, -2, 1) op_1781 (v158[10:0], v447[11:0], v1781[12:0]); // 2.0
    wire [12:0] v1782; shift_adder #(11, 12, 1, 1, 13, 1, 0) op_1782 (v328[10:0], v550[11:0], v1782[12:0]); // 2.0
    wire [12:0] v1783; shift_adder #(11, 12, 1, 1, 13, -1, 0) op_1783 (v264[10:0], v453[11:0], v1783[12:0]); // 2.0
    wire [13:0] v1784; shift_adder #(11, 9, 1, 1, 14, 4, 0) op_1784 (v616[10:0], v538[8:0], v1784[13:0]); // 2.0
    wire [12:0] v1785; shift_adder #(9, 11, 1, 1, 13, -3, 0) op_1785 (v220[8:0], v171[10:0], v1785[12:0]); // 2.0
    wire [10:0] v1786; shift_adder #(9, 9, 1, 1, 11, -1, 0) op_1786 (v575[8:0], v568[8:0], v1786[10:0]); // 2.0
    wire [12:0] v1787; shift_adder #(8, 11, 1, 1, 13, -4, 0) op_1787 (v125[7:0], v145[10:0], v1787[12:0]); // 2.0
    wire [20:0] v1788; shift_adder #(10, 10, 1, 1, 21, -11, 1) op_1788 (v463[9:0], v435[9:0], v1788[20:0]); // 2.0
    wire [20:0] v1789; shift_adder #(12, 19, 1, 1, 21, -9, 0) op_1789 (v434[11:0], v539[18:0], v1789[20:0]); // 2.0
    wire [13:0] v1790; shift_adder #(11, 11, 1, 1, 14, 3, 1) op_1790 (v199[10:0], v169[10:0], v1790[13:0]); // 2.0
    wire [25:0] v1791; shift_adder #(11, 11, 1, 1, 26, 15, 1) op_1791 (v162[10:0], v209[10:0], v1791[25:0]); // 2.0
    wire [18:0] v1792; shift_adder #(18, 11, 1, 1, 19, 7, 0) op_1792 (v493[17:0], v136[10:0], v1792[18:0]); // 2.0
    wire [15:0] v1793; shift_adder #(12, 14, 1, 1, 16, 2, 0) op_1793 (v151[11:0], v481[13:0], v1793[15:0]); // 2.0
    wire [13:0] v1794; shift_adder #(10, 13, 1, 1, 14, -3, 0) op_1794 (v461[9:0], v189[12:0], v1794[13:0]); // 2.0
    wire [15:0] v1795; shift_adder #(13, 12, 1, 1, 16, 4, 0) op_1795 (v346[12:0], v540[11:0], v1795[15:0]); // 2.0
    wire [12:0] v1796; shift_adder #(10, 12, 1, 1, 13, -2, 0) op_1796 (v428[9:0], v224[11:0], v1796[12:0]); // 2.0
    wire [22:0] v1797; shift_adder #(12, 23, 1, 1, 23, -1, 1) op_1797 (v247[11:0], v258[22:0], v1797[22:0]); // 2.0
    wire [22:0] v1798; shift_adder #(22, 12, 1, 1, 23, 10, 0) op_1798 (v617[21:0], v214[11:0], v1798[22:0]); // 2.0
    wire [12:0] v1799; shift_adder #(10, 12, 1, 1, 13, -2, 0) op_1799 (v170[9:0], v553[11:0], v1799[12:0]); // 2.0
    wire [10:0] v1800; shift_adder #(8, 11, 1, 1, 11, 0, 1) op_1800 (v125[7:0], v178[10:0], v1800[10:0]); // 2.0
    wire [18:0] v1801; shift_adder #(11, 11, 1, 1, 19, -8, 1) op_1801 (v241[10:0], v352[10:0], v1801[18:0]); // 2.0
    wire [12:0] v1802; shift_adder #(11, 11, 1, 1, 13, 2, 0) op_1802 (v293[10:0], v131[10:0], v1802[12:0]); // 2.0
    wire [27:0] v1803; shift_adder #(8, 28, 1, 1, 28, -2, 1) op_1803 (v101[7:0], v618[27:0], v1803[27:0]); // 2.0
    wire [16:0] v1804; shift_adder #(8, 17, 1, 1, 17, -8, 1) op_1804 (v119[7:0], v306[16:0], v1804[16:0]); // 2.0
    wire [18:0] v1805; shift_adder #(19, 9, 1, 1, 19, 9, 0) op_1805 (v619[18:0], v620[8:0], v1805[18:0]); // 2.0
    wire [11:0] v1806; shift_adder #(11, 11, 1, 1, 12, 1, 0) op_1806 (v297[10:0], v177[10:0], v1806[11:0]); // 2.0
    wire [23:0] v1807; shift_adder #(11, 11, 1, 1, 24, -13, 1) op_1807 (v144[10:0], v177[10:0], v1807[23:0]); // 2.0
    wire [23:0] v1808; shift_adder #(11, 14, 1, 1, 24, -13, 0) op_1808 (v287[10:0], v290[13:0], v1808[23:0]); // 2.0
    wire [16:0] v1809; shift_adder #(11, 11, 1, 1, 17, 6, 0) op_1809 (v353[10:0], v169[10:0], v1809[16:0]); // 2.0
    wire [10:0] v1810; shift_adder #(8, 11, 1, 1, 11, 0, 1) op_1810 (v105[7:0], v136[10:0], v1810[10:0]); // 2.0
    wire [12:0] v1811; shift_adder #(12, 11, 1, 1, 13, 1, 0) op_1811 (v507[11:0], v213[10:0], v1811[12:0]); // 2.0
    wire [14:0] v1812; shift_adder #(12, 11, 1, 1, 15, -3, 1) op_1812 (v292[11:0], v277[10:0], v1812[14:0]); // 2.0
    wire [13:0] v1813; shift_adder #(11, 12, 1, 1, 14, 2, 1) op_1813 (v197[10:0], v404[11:0], v1813[13:0]); // 2.0
    wire [18:0] v1814; shift_adder #(12, 9, 1, 1, 19, 9, 1) op_1814 (v202[11:0], v370[8:0], v1814[18:0]); // 2.0
    wire [31:0] v1815; shift_adder #(11, 12, 1, 1, 32, 20, 0) op_1815 (v259[10:0], v363[11:0], v1815[31:0]); // 2.0
    wire [15:0] v1816; shift_adder #(12, 12, 1, 1, 16, 4, 0) op_1816 (v382[11:0], v184[11:0], v1816[15:0]); // 2.0
    wire [13:0] v1817; shift_adder #(11, 11, 1, 1, 14, -3, 1) op_1817 (v172[10:0], v518[10:0], v1817[13:0]); // 2.0
    wire [13:0] v1818; shift_adder #(11, 11, 1, 1, 14, 3, 0) op_1818 (v148[10:0], v242[10:0], v1818[13:0]); // 2.0
    wire [12:0] v1819; shift_adder #(11, 12, 1, 1, 13, -1, 1) op_1819 (v328[10:0], v453[11:0], v1819[12:0]); // 2.0
    wire [17:0] v1820; shift_adder #(9, 17, 1, 1, 18, -7, 0) op_1820 (v621[8:0], v545[16:0], v1820[17:0]); // 2.0
    wire [11:0] v1821; shift_adder #(11, 9, 1, 1, 12, 1, 0) op_1821 (v169[10:0], v138[8:0], v1821[11:0]); // 2.0
    wire [11:0] v1822; shift_adder #(11, 10, 1, 1, 12, 1, 0) op_1822 (v622[10:0], v609[9:0], v1822[11:0]); // 2.0
    wire [20:0] v1823; shift_adder #(8, 9, 1, 1, 21, 12, 1) op_1823 (v98[7:0], v351[8:0], v1823[20:0]); // 2.0
    wire [19:0] v1824; shift_adder #(14, 12, 1, 1, 20, -6, 1) op_1824 (v236[13:0], v180[11:0], v1824[19:0]); // 2.0
    wire [12:0] v1825; shift_adder #(11, 11, 1, 1, 13, -2, 0) op_1825 (v418[10:0], v176[10:0], v1825[12:0]); // 2.0
    wire [18:0] v1826; shift_adder #(11, 11, 1, 1, 19, -8, 1) op_1826 (v145[10:0], v393[10:0], v1826[18:0]); // 2.0
    wire [15:0] v1827; shift_adder #(11, 11, 1, 1, 16, 5, 0) op_1827 (v181[10:0], v193[10:0], v1827[15:0]); // 2.0
    wire [14:0] v1828; shift_adder #(12, 12, 1, 1, 15, -3, 0) op_1828 (v383[11:0], v347[11:0], v1828[14:0]); // 2.0
    wire [11:0] v1829; shift_adder #(8, 11, 1, 1, 12, -2, 0) op_1829 (v72[7:0], v191[10:0], v1829[11:0]); // 2.0
    wire [18:0] v1830; shift_adder #(11, 11, 1, 1, 19, -8, 0) op_1830 (v157[10:0], v147[10:0], v1830[18:0]); // 2.0
    wire [15:0] v1831; shift_adder #(11, 14, 1, 1, 16, -5, 0) op_1831 (v602[10:0], v481[13:0], v1831[15:0]); // 2.0
    wire [14:0] v1832; shift_adder #(11, 11, 1, 1, 15, -4, 1) op_1832 (v275[10:0], v301[10:0], v1832[14:0]); // 2.0
    wire [14:0] v1833; shift_adder #(11, 11, 1, 1, 15, -4, 0) op_1833 (v165[10:0], v300[10:0], v1833[14:0]); // 2.0
    wire [13:0] v1834; shift_adder #(11, 11, 1, 1, 14, -3, 1) op_1834 (v195[10:0], v268[10:0], v1834[13:0]); // 2.0
    wire [17:0] v1835; shift_adder #(11, 14, 1, 1, 18, -7, 1) op_1835 (v179[10:0], v481[13:0], v1835[17:0]); // 2.0
    wire [11:0] v1836; shift_adder #(11, 12, 1, 1, 12, 0, 0) op_1836 (v300[10:0], v247[11:0], v1836[11:0]); // 2.0
    wire [23:0] v1837; shift_adder #(11, 22, 1, 1, 24, -13, 0) op_1837 (v131[10:0], v623[21:0], v1837[23:0]); // 2.0
    wire [25:0] v1838; shift_adder #(11, 11, 1, 1, 26, 15, 0) op_1838 (v338[10:0], v168[10:0], v1838[25:0]); // 2.0
    wire [23:0] v1839; shift_adder #(8, 11, 1, 1, 24, -15, 1) op_1839 (v68[7:0], v158[10:0], v1839[23:0]); // 2.0
    wire [15:0] v1840; shift_adder #(11, 11, 1, 1, 16, -5, 0) op_1840 (v209[10:0], v193[10:0], v1840[15:0]); // 2.0
    wire [17:0] v1841; shift_adder #(8, 11, 1, 1, 18, -9, 1) op_1841 (v124[7:0], v303[10:0], v1841[17:0]); // 2.0
    wire [22:0] v1842; shift_adder #(11, 11, 1, 1, 23, 12, 1) op_1842 (v140[10:0], v317[10:0], v1842[22:0]); // 2.0
    wire [21:0] v1843; shift_adder #(21, 13, 1, 1, 22, 9, 0) op_1843 (v624[20:0], v625[12:0], v1843[21:0]); // 2.0
    wire [19:0] v1844; shift_adder #(8, 11, 1, 1, 20, 9, 0) op_1844 (v119[7:0], v287[10:0], v1844[19:0]); // 2.0
    wire [25:0] v1845; shift_adder #(8, 26, 1, 1, 26, -5, 1) op_1845 (v122[7:0], v373[25:0], v1845[25:0]); // 2.0
    wire [17:0] v1846; shift_adder #(11, 14, 1, 1, 18, -7, 0) op_1846 (v190[10:0], v590[13:0], v1846[17:0]); // 2.0
    wire [16:0] v1847; shift_adder #(11, 17, 1, 1, 17, -4, 0) op_1847 (v153[10:0], v615[16:0], v1847[16:0]); // 2.0
    wire [18:0] v1848; shift_adder #(11, 11, 1, 1, 19, -8, 0) op_1848 (v217[10:0], v197[10:0], v1848[18:0]); // 2.0
    wire [14:0] v1849; shift_adder #(10, 11, 1, 1, 15, 4, 0) op_1849 (v626[9:0], v161[10:0], v1849[14:0]); // 2.0
    wire [11:0] v1850; shift_adder #(9, 10, 1, 1, 12, 2, 1) op_1850 (v405[8:0], v222[9:0], v1850[11:0]); // 2.0
    wire [17:0] v1851; shift_adder #(9, 13, 1, 1, 18, -8, 0) op_1851 (v627[8:0], v391[12:0], v1851[17:0]); // 2.0
    wire [11:0] v1852; shift_adder #(11, 11, 1, 1, 12, 1, 0) op_1852 (v375[10:0], v228[10:0], v1852[11:0]); // 2.0
    wire [12:0] v1853; shift_adder #(8, 12, 1, 1, 13, -4, 0) op_1853 (v88[7:0], v434[11:0], v1853[12:0]); // 2.0
    wire [26:0] v1854; shift_adder #(26, 11, 1, 1, 27, 15, 0) op_1854 (v530[25:0], v334[10:0], v1854[26:0]); // 2.0
    wire [21:0] v1855; shift_adder #(8, 13, 1, 1, 22, -13, 1) op_1855 (v126[7:0], v149[12:0], v1855[21:0]); // 2.0
    wire [11:0] v1856; shift_adder #(10, 11, 1, 1, 12, -1, 0) op_1856 (v565[9:0], v297[10:0], v1856[11:0]); // 2.0
    wire [22:0] v1857; shift_adder #(20, 23, 1, 1, 23, -2, 0) op_1857 (v628[19:0], v440[22:0], v1857[22:0]); // 2.0
    wire [14:0] v1858; shift_adder #(11, 11, 1, 1, 15, 4, 1) op_1858 (v238[10:0], v168[10:0], v1858[14:0]); // 2.0
    wire [13:0] v1859; shift_adder #(11, 12, 1, 1, 14, -3, 1) op_1859 (v270[10:0], v382[11:0], v1859[13:0]); // 2.0
    wire [19:0] v1860; shift_adder #(12, 11, 1, 1, 20, 9, 0) op_1860 (v204[11:0], v338[10:0], v1860[19:0]); // 2.0
    wire [14:0] v1861; shift_adder #(12, 12, 1, 1, 15, 3, 1) op_1861 (v321[11:0], v224[11:0], v1861[14:0]); // 2.0
    wire [11:0] v1862; shift_adder #(8, 11, 1, 1, 12, 1, 0) op_1862 (v100[7:0], v234[10:0], v1862[11:0]); // 2.0
    wire [12:0] v1863; shift_adder #(10, 12, 1, 1, 13, -2, 0) op_1863 (v548[9:0], v629[11:0], v1863[12:0]); // 2.0
    wire [20:0] v1864; shift_adder #(11, 12, 1, 1, 21, 9, 0) op_1864 (v297[10:0], v146[11:0], v1864[20:0]); // 2.0
    wire [11:0] v1865; shift_adder #(11, 12, 1, 1, 12, 0, 1) op_1865 (v131[10:0], v285[11:0], v1865[11:0]); // 2.0
    wire [11:0] v1866; shift_adder #(11, 10, 1, 1, 12, 1, 0) op_1866 (v324[10:0], v501[9:0], v1866[11:0]); // 2.0
    wire [14:0] v1867; shift_adder #(11, 12, 1, 1, 15, 3, 1) op_1867 (v178[10:0], v553[11:0], v1867[14:0]); // 2.0
    wire [10:0] v1868; shift_adder #(11, 9, 1, 1, 11, 0, 0) op_1868 (v244[10:0], v561[8:0], v1868[10:0]); // 2.0
    wire [17:0] v1869; shift_adder #(8, 15, 1, 1, 18, 3, 0) op_1869 (v98[7:0], v630[14:0], v1869[17:0]); // 2.0
    wire [33:0] v1870; shift_adder #(13, 10, 1, 1, 34, -21, 1) op_1870 (v631[12:0], v527[9:0], v1870[33:0]); // 2.0
    wire [11:0] v1871; shift_adder #(10, 11, 1, 1, 12, -1, 0) op_1871 (v445[9:0], v229[10:0], v1871[11:0]); // 2.0
    wire [12:0] v1872; shift_adder #(11, 12, 1, 1, 13, -2, 0) op_1872 (v329[10:0], v207[11:0], v1872[12:0]); // 2.0
    wire [11:0] v1873; shift_adder #(12, 11, 1, 1, 12, 0, 0) op_1873 (v227[11:0], v136[10:0], v1873[11:0]); // 2.0
    wire [14:0] v1874; shift_adder #(8, 14, 1, 1, 15, -6, 0) op_1874 (v87[7:0], v412[13:0], v1874[14:0]); // 2.0
    wire [24:0] v1875; shift_adder #(8, 25, 1, 1, 25, -10, 0) op_1875 (v84[7:0], v611[24:0], v1875[24:0]); // 2.0
    wire [32:0] v1876; shift_adder #(8, 12, 1, 1, 33, 21, 1) op_1876 (v108[7:0], v365[11:0], v1876[32:0]); // 2.0
    wire [10:0] v1877; shift_adder #(9, 10, 1, 1, 11, -1, 0) op_1877 (v503[8:0], v606[9:0], v1877[10:0]); // 2.0
    wire [26:0] v1878; shift_adder #(11, 11, 1, 1, 27, -16, 1) op_1878 (v294[10:0], v139[10:0], v1878[26:0]); // 2.0
    wire [14:0] v1879; shift_adder #(11, 11, 1, 1, 15, -4, 1) op_1879 (v232[10:0], v197[10:0], v1879[14:0]); // 2.0
    wire [14:0] v1880; shift_adder #(8, 9, 1, 1, 15, 5, 1) op_1880 (v81[7:0], v351[8:0], v1880[14:0]); // 2.0
    wire [25:0] v1881; shift_adder #(11, 11, 1, 1, 26, 15, 1) op_1881 (v131[10:0], v178[10:0], v1881[25:0]); // 2.0
    wire [25:0] v1882; shift_adder #(11, 18, 1, 1, 26, -15, 1) op_1882 (v323[10:0], v633[17:0], v1882[25:0]); // 2.0
    wire [16:0] v1883; shift_adder #(11, 16, 1, 1, 17, -6, 0) op_1883 (v148[10:0], v634[15:0], v1883[16:0]); // 2.0
    wire [17:0] v1884; shift_adder #(8, 18, 1, 1, 18, 0, 1) op_1884 (v80[7:0], v494[17:0], v1884[17:0]); // 2.0
    wire [21:0] v1885; shift_adder #(8, 11, 1, 1, 22, 11, 0) op_1885 (v112[7:0], v145[10:0], v1885[21:0]); // 2.0
    wire [19:0] v1886; shift_adder #(11, 15, 1, 1, 20, 5, 1) op_1886 (v187[10:0], v318[14:0], v1886[19:0]); // 2.0
    wire [15:0] v1887; shift_adder #(14, 11, 1, 1, 16, -2, 0) op_1887 (v555[13:0], v152[10:0], v1887[15:0]); // 2.0
    wire [11:0] v1888; shift_adder #(11, 11, 1, 1, 12, 0, 1) op_1888 (v211[10:0], v379[10:0], v1888[11:0]); // 2.0
    wire [15:0] v1889; shift_adder #(11, 11, 1, 1, 16, -5, 1) op_1889 (v216[10:0], v199[10:0], v1889[15:0]); // 2.0
    wire [17:0] v1890; shift_adder #(8, 11, 1, 1, 18, -9, 1) op_1890 (v123[7:0], v338[10:0], v1890[17:0]); // 2.0
    wire [13:0] v1891; shift_adder #(12, 10, 1, 1, 14, 3, 0) op_1891 (v285[11:0], v509[9:0], v1891[13:0]); // 2.0
    wire [12:0] v1892; shift_adder #(11, 13, 1, 1, 13, -1, 0) op_1892 (v142[10:0], v406[12:0], v1892[12:0]); // 2.0
    wire [11:0] v1893; shift_adder #(11, 11, 1, 1, 12, 1, 1) op_1893 (v172[10:0], v303[10:0], v1893[11:0]); // 2.0
    wire [10:0] v1894; shift_adder #(11, 10, 1, 1, 11, 0, 0) op_1894 (v455[10:0], v463[9:0], v1894[10:0]); // 2.0
    wire [20:0] v1895; shift_adder #(12, 12, 1, 1, 21, 9, 0) op_1895 (v137[11:0], v304[11:0], v1895[20:0]); // 2.0
    wire [31:0] v1896; shift_adder #(11, 30, 1, 1, 32, 2, 0) op_1896 (v241[10:0], v605[29:0], v1896[31:0]); // 2.0
    wire [15:0] v1897; shift_adder #(11, 11, 1, 1, 16, 5, 0) op_1897 (v259[10:0], v379[10:0], v1897[15:0]); // 2.0
    wire [11:0] v1898; shift_adder #(11, 11, 1, 1, 12, 1, 0) op_1898 (v396[10:0], v206[10:0], v1898[11:0]); // 2.0
    wire [15:0] v1899; shift_adder #(11, 11, 1, 1, 16, 5, 0) op_1899 (v195[10:0], v361[10:0], v1899[15:0]); // 2.0
    wire [18:0] v1900; shift_adder #(11, 9, 1, 1, 19, 9, 0) op_1900 (v245[10:0], v138[8:0], v1900[18:0]); // 2.0
    wire [12:0] v1901; shift_adder #(11, 11, 1, 1, 13, 2, 0) op_1901 (v178[10:0], v150[10:0], v1901[12:0]); // 2.0
    wire [19:0] v1902; shift_adder #(8, 12, 1, 1, 20, 8, 0) op_1902 (v117[7:0], v552[11:0], v1902[19:0]); // 2.0
    wire [22:0] v1903; shift_adder #(23, 10, 1, 1, 23, 12, 0) op_1903 (v635[22:0], v260[9:0], v1903[22:0]); // 2.0
    wire [14:0] v1904; shift_adder #(11, 11, 1, 1, 15, 4, 1) op_1904 (v157[10:0], v219[10:0], v1904[14:0]); // 2.0
    wire [10:0] v1905; shift_adder #(8, 11, 1, 1, 11, 0, 0) op_1905 (v108[7:0], v415[10:0], v1905[10:0]); // 2.0
    wire [11:0] v1906; shift_adder #(11, 11, 1, 1, 12, 1, 0) op_1906 (v244[10:0], v283[10:0], v1906[11:0]); // 2.0
    wire [12:0] v1907; shift_adder #(11, 10, 1, 1, 13, -2, 0) op_1907 (v362[10:0], v235[9:0], v1907[12:0]); // 2.0
    wire [12:0] v1908; shift_adder #(11, 10, 1, 1, 13, 3, 0) op_1908 (v297[10:0], v554[9:0], v1908[12:0]); // 2.0
    wire [12:0] v1909; shift_adder #(12, 9, 1, 1, 13, 3, 0) op_1909 (v457[11:0], v637[8:0], v1909[12:0]); // 2.0
    wire [16:0] v1910; shift_adder #(11, 15, 1, 1, 17, -6, 0) op_1910 (v229[10:0], v456[14:0], v1910[16:0]); // 2.0
    wire [12:0] v1911; shift_adder #(9, 11, 1, 1, 13, -3, 0) op_1911 (v395[8:0], v600[10:0], v1911[12:0]); // 2.0
    wire [15:0] v1912; shift_adder #(14, 12, 1, 1, 16, 4, 0) op_1912 (v638[13:0], v457[11:0], v1912[15:0]); // 2.0
    wire [15:0] v1913; shift_adder #(11, 11, 1, 1, 16, 5, 0) op_1913 (v155[10:0], v136[10:0], v1913[15:0]); // 2.0
    wire [12:0] v1914; shift_adder #(10, 10, 1, 1, 13, -3, 0) op_1914 (v421[9:0], v282[9:0], v1914[12:0]); // 2.0
    wire [11:0] v1915; shift_adder #(10, 12, 1, 1, 12, 0, 0) op_1915 (v639[9:0], v292[11:0], v1915[11:0]); // 2.0
    wire [12:0] v1916; shift_adder #(10, 12, 1, 1, 13, -2, 0) op_1916 (v421[9:0], v589[11:0], v1916[12:0]); // 2.0
    wire [18:0] v1917; shift_adder #(9, 19, 1, 1, 19, -8, 0) op_1917 (v230[8:0], v640[18:0], v1917[18:0]); // 2.0
    wire [33:0] v1918; shift_adder #(31, 33, 1, 1, 34, -3, 0) op_1918 (v641[30:0], v608[32:0], v1918[33:0]); // 2.0
    wire [14:0] v1919; shift_adder #(11, 11, 1, 1, 15, 4, 0) op_1919 (v270[10:0], v215[10:0], v1919[14:0]); // 2.0
    wire [15:0] v1920; shift_adder #(16, 11, 1, 1, 16, 2, 0) op_1920 (v504[15:0], v232[10:0], v1920[15:0]); // 2.0
    wire [14:0] v1921; shift_adder #(14, 12, 1, 1, 15, -1, 0) op_1921 (v460[13:0], v642[11:0], v1921[14:0]); // 2.0
    wire [11:0] v1922; shift_adder #(11, 11, 1, 1, 12, 0, 0) op_1922 (v320[10:0], v158[10:0], v1922[11:0]); // 2.0
    wire [11:0] v1923; shift_adder #(8, 11, 1, 1, 12, 1, 0) op_1923 (v116[7:0], v241[10:0], v1923[11:0]); // 2.0
    wire [12:0] v1924; shift_adder #(11, 12, 1, 1, 13, 1, 0) op_1924 (v132[10:0], v164[11:0], v1924[12:0]); // 2.0
    wire [24:0] v1925; shift_adder #(14, 18, 1, 1, 25, 7, 0) op_1925 (v290[13:0], v633[17:0], v1925[24:0]); // 2.0
    wire [20:0] v1926; shift_adder #(12, 10, 1, 1, 21, -9, 0) op_1926 (v473[11:0], v643[9:0], v1926[20:0]); // 2.0
    wire [13:0] v1927; shift_adder #(11, 11, 1, 1, 14, -3, 1) op_1927 (v268[10:0], v187[10:0], v1927[13:0]); // 2.0
    wire [15:0] v1928; shift_adder #(11, 14, 1, 1, 16, -5, 0) op_1928 (v131[10:0], v410[13:0], v1928[15:0]); // 2.0
    wire [15:0] v1929; shift_adder #(11, 16, 1, 1, 16, -4, 0) op_1929 (v195[10:0], v519[15:0], v1929[15:0]); // 2.0
    wire [22:0] v1930; shift_adder #(11, 12, 1, 1, 23, 11, 0) op_1930 (v195[10:0], v447[11:0], v1930[22:0]); // 2.0
    wire [18:0] v1931; shift_adder #(11, 19, 1, 1, 19, -7, 0) op_1931 (v345[10:0], v558[18:0], v1931[18:0]); // 2.0
    wire [14:0] v1932; shift_adder #(11, 12, 1, 1, 15, 3, 1) op_1932 (v188[10:0], v409[11:0], v1932[14:0]); // 2.0
    wire [14:0] v1933; shift_adder #(15, 13, 1, 1, 15, 0, 0) op_1933 (v253[14:0], v645[12:0], v1933[14:0]); // 2.0
    wire [13:0] v1934; shift_adder #(12, 13, 1, 1, 14, -1, 0) op_1934 (v151[11:0], v391[12:0], v1934[13:0]); // 2.0
    wire [24:0] v1935; shift_adder #(8, 11, 1, 1, 25, -16, 1) op_1935 (v92[7:0], v238[10:0], v1935[24:0]); // 2.0
    wire [22:0] v1936; shift_adder #(11, 23, 1, 1, 23, -10, 0) op_1936 (v241[10:0], v564[22:0], v1936[22:0]); // 2.0
    wire [16:0] v1937; shift_adder #(11, 11, 1, 1, 17, -6, 1) op_1937 (v289[10:0], v153[10:0], v1937[16:0]); // 2.0
    wire [17:0] v1938; shift_adder #(10, 18, 1, 1, 18, -7, 0) op_1938 (v366[9:0], v535[17:0], v1938[17:0]); // 2.0
    wire [13:0] v1939; shift_adder #(11, 11, 1, 1, 14, -3, 0) op_1939 (v293[10:0], v197[10:0], v1939[13:0]); // 2.0
    wire [11:0] v1940; shift_adder #(8, 10, 1, 1, 12, -3, 0) op_1940 (v105[7:0], v311[9:0], v1940[11:0]); // 2.0
    wire [12:0] v1941; shift_adder #(11, 11, 1, 1, 13, 2, 1) op_1941 (v250[10:0], v352[10:0], v1941[12:0]); // 2.0
    wire [18:0] v1942; shift_adder #(8, 12, 1, 1, 19, -10, 1) op_1942 (v120[7:0], v423[11:0], v1942[18:0]); // 2.0
    wire [10:0] v1943; shift_adder #(8, 11, 1, 1, 11, -1, 0) op_1943 (v98[7:0], v233[10:0], v1943[10:0]); // 2.0
    wire [13:0] v1944; shift_adder #(12, 13, 1, 1, 14, 1, 0) op_1944 (v321[11:0], v625[12:0], v1944[13:0]); // 2.0
    wire [18:0] v1945; shift_adder #(11, 11, 1, 1, 19, 8, 0) op_1945 (v375[10:0], v187[10:0], v1945[18:0]); // 2.0
    wire [12:0] v1946; shift_adder #(11, 12, 1, 1, 13, -1, 0) op_1946 (v165[10:0], v397[11:0], v1946[12:0]); // 2.0
    wire [14:0] v1947; shift_adder #(11, 15, 1, 1, 15, -3, 1) op_1947 (v269[10:0], v318[14:0], v1947[14:0]); // 2.0
    wire [11:0] v1948; shift_adder #(9, 11, 1, 1, 12, 1, 0) op_1948 (v627[8:0], v148[10:0], v1948[11:0]); // 2.0
    wire [12:0] v1949; shift_adder #(8, 13, 1, 1, 13, -3, 1) op_1949 (v81[7:0], v272[12:0], v1949[12:0]); // 2.0
    wire [15:0] v1950; shift_adder #(16, 11, 1, 1, 16, 3, 0) op_1950 (v166[15:0], v644[10:0], v1950[15:0]); // 2.0
    wire [11:0] v1951; shift_adder #(9, 12, 1, 1, 12, -1, 0) op_1951 (v405[8:0], v146[11:0], v1951[11:0]); // 2.0
    wire [28:0] v1952; shift_adder #(12, 12, 1, 1, 29, 17, 1) op_1952 (v380[11:0], v582[11:0], v1952[28:0]); // 2.0
    wire [32:0] v1953; shift_adder #(11, 10, 1, 1, 33, 23, 0) op_1953 (v251[10:0], v450[9:0], v1953[32:0]); // 2.0
    wire [22:0] v1954; shift_adder #(8, 11, 1, 1, 23, -14, 1) op_1954 (v104[7:0], v425[10:0], v1954[22:0]); // 2.0
    wire [12:0] v1955; shift_adder #(13, 11, 1, 1, 13, 1, 0) op_1955 (v646[12:0], v175[10:0], v1955[12:0]); // 2.0
    wire [11:0] v1956; shift_adder #(10, 10, 1, 1, 12, 1, 0) op_1956 (v647[9:0], v648[9:0], v1956[11:0]); // 2.0
    wire [11:0] v1957; shift_adder #(10, 9, 1, 1, 12, 2, 0) op_1957 (v225[9:0], v508[8:0], v1957[11:0]); // 2.0
    wire [11:0] v1958; shift_adder #(11, 11, 1, 1, 12, 0, 0) op_1958 (v188[10:0], v129[10:0], v1958[11:0]); // 2.0
    wire [35:0] v1959; shift_adder #(15, 12, 1, 1, 36, -21, 1) op_1959 (v649[14:0], v650[11:0], v1959[35:0]); // 2.0
    wire [10:0] v1960; shift_adder #(11, 9, 1, 1, 11, 0, 0) op_1960 (v203[10:0], v651[8:0], v1960[10:0]); // 2.0
    wire [15:0] v1961; shift_adder #(9, 15, 1, 1, 16, -6, 0) op_1961 (v302[8:0], v652[14:0], v1961[15:0]); // 2.0
    wire [13:0] v1962; shift_adder #(11, 12, 1, 1, 14, -3, 0) op_1962 (v274[10:0], v336[11:0], v1962[13:0]); // 2.0
    wire [11:0] v1963; shift_adder #(11, 12, 1, 1, 12, 0, 0) op_1963 (v312[10:0], v339[11:0], v1963[11:0]); // 2.0
    wire [14:0] v1964; shift_adder #(11, 11, 1, 1, 15, 4, 1) op_1964 (v294[10:0], v375[10:0], v1964[14:0]); // 2.0
    wire [10:0] v1965; shift_adder #(10, 11, 1, 1, 11, 0, 0) op_1965 (v435[9:0], v187[10:0], v1965[10:0]); // 2.0
    wire [18:0] v1966; shift_adder #(11, 11, 1, 1, 19, -8, 0) op_1966 (v203[10:0], v162[10:0], v1966[18:0]); // 2.0
    wire [12:0] v1967; shift_adder #(12, 11, 1, 1, 13, 2, 0) op_1967 (v452[11:0], v653[10:0], v1967[12:0]); // 2.0
    wire [12:0] v1968; shift_adder #(10, 11, 1, 1, 13, -3, 0) op_1968 (v263[9:0], v245[10:0], v1968[12:0]); // 2.0
    wire [15:0] v1969; shift_adder #(13, 16, 1, 1, 16, -2, 0) op_1969 (v654[12:0], v655[15:0], v1969[15:0]); // 2.0
    wire [12:0] v1970; shift_adder #(10, 11, 1, 1, 13, -2, 0) op_1970 (v446[9:0], v424[10:0], v1970[12:0]); // 2.0
    wire [22:0] v1971; shift_adder #(22, 9, 1, 1, 23, 13, 0) op_1971 (v656[21:0], v531[8:0], v1971[22:0]); // 2.0
    wire [13:0] v1972; shift_adder #(11, 12, 1, 1, 14, -3, 0) op_1972 (v141[10:0], v523[11:0], v1972[13:0]); // 2.0
    wire [13:0] v1973; shift_adder #(8, 11, 1, 1, 14, -5, 0) op_1973 (v100[7:0], v317[10:0], v1973[13:0]); // 2.0
    wire [12:0] v1974; shift_adder #(12, 12, 1, 1, 13, 0, 0) op_1974 (v657[11:0], v194[11:0], v1974[12:0]); // 2.0
    wire [14:0] v1975; shift_adder #(9, 14, 1, 1, 15, -5, 0) op_1975 (v322[8:0], v658[13:0], v1975[14:0]); // 2.0
    wire [20:0] v1976; shift_adder #(11, 11, 1, 1, 21, -10, 1) op_1976 (v264[10:0], v217[10:0], v1976[20:0]); // 2.0
    wire [11:0] v1977; shift_adder #(8, 11, 1, 1, 12, -3, 1) op_1977 (v69[7:0], v352[10:0], v1977[11:0]); // 2.0
    wire [17:0] v1978; shift_adder #(8, 11, 1, 1, 18, 7, 0) op_1978 (v102[7:0], v319[10:0], v1978[17:0]); // 2.0
    wire [13:0] v1979; shift_adder #(10, 12, 1, 1, 14, -4, 0) op_1979 (v606[9:0], v382[11:0], v1979[13:0]); // 2.0
    wire [13:0] v1980; shift_adder #(11, 13, 1, 1, 14, -3, 0) op_1980 (v188[10:0], v458[12:0], v1980[13:0]); // 2.0
    wire [20:0] v1981; shift_adder #(11, 11, 1, 1, 21, 10, 1) op_1981 (v162[10:0], v233[10:0], v1981[20:0]); // 2.0
    wire [13:0] v1982; shift_adder #(11, 12, 1, 1, 14, -3, 0) op_1982 (v156[10:0], v540[11:0], v1982[13:0]); // 2.0
    wire [19:0] v1983; shift_adder #(8, 15, 1, 1, 20, 5, 1) op_1983 (v104[7:0], v528[14:0], v1983[19:0]); // 2.0
    wire [19:0] v1984; shift_adder #(11, 11, 1, 1, 20, 9, 1) op_1984 (v374[10:0], v324[10:0], v1984[19:0]); // 2.0
    wire [12:0] v1985; shift_adder #(13, 10, 1, 1, 13, 2, 0) op_1985 (v476[12:0], v428[9:0], v1985[12:0]); // 2.0
    wire [11:0] v1986; shift_adder #(11, 12, 1, 1, 12, 0, 1) op_1986 (v233[10:0], v434[11:0], v1986[11:0]); // 2.0
    wire [17:0] v1987; shift_adder #(11, 11, 1, 1, 18, 7, 1) op_1987 (v147[10:0], v139[10:0], v1987[17:0]); // 2.0
    wire [21:0] v1988; shift_adder #(11, 9, 1, 1, 22, 13, 1) op_1988 (v251[10:0], v370[8:0], v1988[21:0]); // 2.0
    wire [26:0] v1989; shift_adder #(11, 12, 1, 1, 27, 15, 0) op_1989 (v131[10:0], v553[11:0], v1989[26:0]); // 2.0
    wire [11:0] v1990; shift_adder #(11, 11, 1, 1, 12, 0, 0) op_1990 (v418[10:0], v277[10:0], v1990[11:0]); // 2.0
    wire [16:0] v1991; shift_adder #(14, 17, 1, 1, 17, -2, 0) op_1991 (v236[13:0], v306[16:0], v1991[16:0]); // 2.0
    wire [12:0] v1992; shift_adder #(12, 11, 1, 1, 13, 1, 0) op_1992 (v180[11:0], v317[10:0], v1992[12:0]); // 2.0
    wire [22:0] v1993; shift_adder #(12, 12, 1, 1, 23, -11, 1) op_1993 (v550[11:0], v447[11:0], v1993[22:0]); // 2.0
    wire [28:0] v1994; shift_adder #(28, 13, 1, 1, 29, 15, 0) op_1994 (v618[27:0], v660[12:0], v1994[28:0]); // 2.0
    wire [11:0] v1995; shift_adder #(12, 11, 1, 1, 12, 0, 0) op_1995 (v363[11:0], v237[10:0], v1995[11:0]); // 2.0
    wire [11:0] v1996; shift_adder #(9, 11, 1, 1, 12, 1, 0) op_1996 (v231[8:0], v602[10:0], v1996[11:0]); // 2.0
    wire [12:0] v1997; shift_adder #(10, 11, 1, 1, 13, -2, 0) op_1997 (v548[9:0], v276[10:0], v1997[12:0]); // 2.0
    wire [12:0] v1998; shift_adder #(11, 12, 1, 1, 13, -1, 0) op_1998 (v200[10:0], v363[11:0], v1998[12:0]); // 2.0
    wire [18:0] v1999; shift_adder #(10, 18, 1, 1, 19, -8, 0) op_1999 (v606[9:0], v286[17:0], v1999[18:0]); // 2.0
    wire [11:0] v2000; shift_adder #(12, 10, 1, 1, 12, 0, 0) op_2000 (v614[11:0], v520[9:0], v2000[11:0]); // 2.0
    wire [11:0] v2001; shift_adder #(11, 11, 1, 1, 12, 0, 0) op_2001 (v661[10:0], v338[10:0], v2001[11:0]); // 2.0
    wire [12:0] v2002; shift_adder #(9, 12, 1, 1, 13, -3, 0) op_2002 (v128[8:0], v137[11:0], v2002[12:0]); // 2.0
    wire [14:0] v2003; shift_adder #(12, 14, 1, 1, 15, -2, 1) op_2003 (v214[11:0], v590[13:0], v2003[14:0]); // 2.0
    wire [11:0] v2004; shift_adder #(9, 11, 1, 1, 12, -2, 0) op_2004 (v340[8:0], v662[10:0], v2004[11:0]); // 2.0
    wire [14:0] v2005; shift_adder #(11, 11, 1, 1, 15, -4, 1) op_2005 (v319[10:0], v328[10:0], v2005[14:0]); // 2.0
    wire [23:0] v2006; shift_adder #(11, 22, 1, 1, 24, -13, 0) op_2006 (v455[10:0], v371[21:0], v2006[23:0]); // 2.0
    wire [16:0] v2007; shift_adder #(9, 16, 1, 1, 17, -7, 0) op_2007 (v663[8:0], v566[15:0], v2007[16:0]); // 2.0
    wire [13:0] v2008; shift_adder #(11, 11, 1, 1, 14, -3, 0) op_2008 (v210[10:0], v320[10:0], v2008[13:0]); // 2.0
    wire [24:0] v2009; shift_adder #(8, 11, 1, 1, 25, 14, 1) op_2009 (v68[7:0], v190[10:0], v2009[24:0]); // 2.0
    wire [12:0] v2010; shift_adder #(11, 13, 1, 1, 13, 0, 0) op_2010 (v191[10:0], v189[12:0], v2010[12:0]); // 2.0
    wire [13:0] v2011; shift_adder #(12, 11, 1, 1, 14, 3, 0) op_2011 (v457[11:0], v154[10:0], v2011[13:0]); // 2.0
    wire [29:0] v2012; shift_adder #(9, 8, 1, 1, 30, 21, 1) op_2012 (v405[8:0], v97[7:0], v2012[29:0]); // 2.0
    wire [17:0] v2013; shift_adder #(11, 11, 1, 1, 18, 7, 0) op_2013 (v334[10:0], v134[10:0], v2013[17:0]); // 2.0
    wire [12:0] v2014; shift_adder #(12, 11, 1, 1, 13, 1, 0) op_2014 (v664[11:0], v334[10:0], v2014[12:0]); // 2.0
    wire [14:0] v2015; shift_adder #(12, 14, 1, 1, 15, -2, 1) op_2015 (v550[11:0], v271[13:0], v2015[14:0]); // 2.0
    wire [14:0] v2016; shift_adder #(11, 13, 1, 1, 15, 2, 0) op_2016 (v200[10:0], v406[12:0], v2016[14:0]); // 2.0
    wire [11:0] v2017; shift_adder #(8, 12, 1, 1, 12, -2, 0) op_2017 (v119[7:0], v382[11:0], v2017[11:0]); // 2.0
    wire [12:0] v2018; shift_adder #(12, 11, 1, 1, 13, 1, 0) op_2018 (v657[11:0], v317[10:0], v2018[12:0]); // 2.0
    wire [11:0] v2019; shift_adder #(8, 11, 1, 1, 12, -2, 0) op_2019 (v127[7:0], v283[10:0], v2019[11:0]); // 2.0
    wire [14:0] v2020; shift_adder #(14, 11, 1, 1, 15, 4, 0) op_2020 (v665[13:0], v155[10:0], v2020[14:0]); // 2.0
    wire [18:0] v2021; shift_adder #(17, 12, 1, 1, 19, 7, 0) op_2021 (v414[16:0], v397[11:0], v2021[18:0]); // 2.0
    wire [14:0] v2022; shift_adder #(11, 11, 1, 1, 15, -4, 0) op_2022 (v210[10:0], v153[10:0], v2022[14:0]); // 2.0
    wire [21:0] v2023; shift_adder #(11, 11, 1, 1, 22, 11, 1) op_2023 (v396[10:0], v367[10:0], v2023[21:0]); // 2.0
    wire [12:0] v2024; shift_adder #(10, 12, 1, 1, 13, 1, 0) op_2024 (v666[9:0], v383[11:0], v2024[12:0]); // 2.0
    wire [17:0] v2025; shift_adder #(11, 12, 1, 1, 18, 6, 0) op_2025 (v136[10:0], v292[11:0], v2025[17:0]); // 2.0
    wire [24:0] v2026; shift_adder #(11, 11, 1, 1, 25, 14, 0) op_2026 (v171[10:0], v135[10:0], v2026[24:0]); // 2.0
    wire [11:0] v2027; shift_adder #(11, 11, 1, 1, 12, -1, 0) op_2027 (v250[10:0], v182[10:0], v2027[11:0]); // 2.0
    wire [13:0] v2028; shift_adder #(12, 11, 1, 1, 14, -2, 0) op_2028 (v544[11:0], v213[10:0], v2028[13:0]); // 2.0
    wire [27:0] v2029; shift_adder #(8, 11, 1, 1, 28, -19, 0) op_2029 (v111[7:0], v187[10:0], v2029[27:0]); // 2.0
    wire [11:0] v2030; shift_adder #(12, 11, 1, 1, 12, 0, 0) op_2030 (v347[11:0], v341[10:0], v2030[11:0]); // 2.0
    wire [12:0] v2031; shift_adder #(11, 12, 1, 1, 13, -2, 1) op_2031 (v210[10:0], v500[11:0], v2031[12:0]); // 2.0
    wire [21:0] v2032; shift_adder #(11, 14, 1, 1, 22, 8, 0) op_2032 (v156[10:0], v290[13:0], v2032[21:0]); // 2.0
    wire [11:0] v2033; shift_adder #(11, 11, 1, 1, 12, -1, 1) op_2033 (v241[10:0], v297[10:0], v2033[11:0]); // 2.0
    wire [18:0] v2034; shift_adder #(11, 11, 1, 1, 19, 8, 0) op_2034 (v319[10:0], v293[10:0], v2034[18:0]); // 2.0
    wire [12:0] v2035; shift_adder #(12, 11, 1, 1, 13, 2, 0) op_2035 (v321[11:0], v386[10:0], v2035[12:0]); // 2.0
    wire [13:0] v2036; shift_adder #(12, 13, 1, 1, 14, -1, 0) op_2036 (v183[11:0], v344[12:0], v2036[13:0]); // 2.0
    wire [14:0] v2037; shift_adder #(11, 11, 1, 1, 15, -4, 0) op_2037 (v213[10:0], v379[10:0], v2037[14:0]); // 2.0
    wire [20:0] v2038; shift_adder #(17, 20, 1, 1, 21, -3, 0) op_2038 (v551[16:0], v484[19:0], v2038[20:0]); // 2.0
    wire [11:0] v2039; shift_adder #(11, 10, 1, 1, 12, 1, 1) op_2039 (v156[10:0], v592[9:0], v2039[11:0]); // 2.0
    wire [13:0] v2040; shift_adder #(11, 9, 1, 1, 14, 4, 1) op_2040 (v209[10:0], v302[8:0], v2040[13:0]); // 2.0
    wire [23:0] v2041; shift_adder #(11, 11, 1, 1, 24, 13, 0) op_2041 (v269[10:0], v163[10:0], v2041[23:0]); // 2.0
    wire [21:0] v2042; shift_adder #(22, 17, 1, 1, 22, 4, 0) op_2042 (v656[21:0], v667[16:0], v2042[21:0]); // 2.0
    wire [11:0] v2043; shift_adder #(11, 11, 1, 1, 12, -1, 0) op_2043 (v264[10:0], v275[10:0], v2043[11:0]); // 2.0
    wire [14:0] v2044; shift_adder #(11, 11, 1, 1, 15, 4, 1) op_2044 (v251[10:0], v176[10:0], v2044[14:0]); // 2.0
    wire [13:0] v2045; shift_adder #(12, 12, 1, 1, 14, -2, 0) op_2045 (v579[11:0], v314[11:0], v2045[13:0]); // 2.0
    wire [14:0] v2046; shift_adder #(11, 11, 1, 1, 15, 4, 1) op_2046 (v158[10:0], v206[10:0], v2046[14:0]); // 2.0
    wire [17:0] v2047; shift_adder #(12, 12, 1, 1, 18, -6, 1) op_2047 (v365[11:0], v365[11:0], v2047[17:0]); // 2.0
    wire [13:0] v2048; shift_adder #(12, 12, 1, 1, 14, -2, 1) op_2048 (v257[11:0], v380[11:0], v2048[13:0]); // 2.0
    wire [13:0] v2049; shift_adder #(12, 10, 1, 1, 14, 4, 0) op_2049 (v668[11:0], v291[9:0], v2049[13:0]); // 2.0
    wire [35:0] v2050; shift_adder #(33, 11, 1, 1, 36, 25, 0) op_2050 (v608[32:0], v659[10:0], v2050[35:0]); // 2.0
    wire [10:0] v2051; shift_adder #(9, 11, 1, 1, 11, 0, 0) op_2051 (v221[8:0], v210[10:0], v2051[10:0]); // 2.0
    wire [18:0] v2052; shift_adder #(11, 11, 1, 1, 19, 8, 1) op_2052 (v223[10:0], v182[10:0], v2052[18:0]); // 2.0
    wire [14:0] v2053; shift_adder #(13, 10, 1, 1, 15, 4, 0) op_2053 (v149[12:0], v554[9:0], v2053[14:0]); // 2.0
    wire [10:0] v2054; shift_adder #(10, 11, 1, 1, 11, 0, 0) op_2054 (v260[9:0], v210[10:0], v2054[10:0]); // 2.0
    wire [19:0] v2055; shift_adder #(18, 13, 1, 1, 20, 7, 0) op_2055 (v562[17:0], v326[12:0], v2055[19:0]); // 2.0
    wire [13:0] v2056; shift_adder #(8, 10, 1, 1, 14, -5, 1) op_2056 (v79[7:0], v610[9:0], v2056[13:0]); // 2.0
    wire [34:0] v2057; shift_adder #(10, 35, 1, 1, 35, -24, 0) op_2057 (v669[9:0], v670[34:0], v2057[34:0]); // 2.0
    wire [36:0] v2058; shift_adder #(11, 11, 1, 1, 37, -26, 1) op_2058 (v671[10:0], v396[10:0], v2058[36:0]); // 2.0
    wire [11:0] v2059; shift_adder #(11, 11, 1, 1, 12, -1, 0) op_2059 (v644[10:0], v672[10:0], v2059[11:0]); // 2.0
    wire [14:0] v2060; shift_adder #(12, 13, 1, 1, 15, -3, 0) op_2060 (v174[11:0], v344[12:0], v2060[14:0]); // 2.0
    wire [11:0] v2061; shift_adder #(11, 11, 1, 1, 12, 0, 0) op_2061 (v195[10:0], v132[10:0], v2061[11:0]); // 2.0
    wire [12:0] v2062; shift_adder #(13, 11, 1, 1, 13, 0, 0) op_2062 (v645[12:0], v208[10:0], v2062[12:0]); // 2.0
    wire [11:0] v2063; shift_adder #(11, 11, 1, 1, 12, 0, 0) op_2063 (v219[10:0], v237[10:0], v2063[11:0]); // 2.0
    wire [11:0] v2064; shift_adder #(11, 11, 1, 1, 12, 0, 0) op_2064 (v145[10:0], v600[10:0], v2064[11:0]); // 2.0
    wire [12:0] v2065; shift_adder #(11, 11, 1, 1, 13, 2, 1) op_2065 (v173[10:0], v393[10:0], v2065[12:0]); // 2.0
    wire [12:0] v2066; shift_adder #(11, 11, 1, 1, 13, 2, 0) op_2066 (v289[10:0], v367[10:0], v2066[12:0]); // 2.0
    wire [13:0] v2067; shift_adder #(11, 13, 1, 1, 14, -3, 0) op_2067 (v505[10:0], v189[12:0], v2067[13:0]); // 2.0
    wire [14:0] v2068; shift_adder #(12, 11, 1, 1, 15, -3, 1) op_2068 (v174[11:0], v255[10:0], v2068[14:0]); // 2.0
    wire [16:0] v2069; shift_adder #(11, 11, 1, 1, 17, 6, 0) op_2069 (v334[10:0], v264[10:0], v2069[16:0]); // 2.0
    wire [20:0] v2070; shift_adder #(19, 19, 1, 1, 21, -2, 0) op_2070 (v558[18:0], v597[18:0], v2070[20:0]); // 2.0
    wire [11:0] v2071; shift_adder #(11, 11, 1, 1, 12, 0, 1) op_2071 (v158[10:0], v132[10:0], v2071[11:0]); // 2.0
    wire [11:0] v2072; shift_adder #(8, 10, 1, 1, 12, 2, 0) op_2072 (v105[7:0], v366[9:0], v2072[11:0]); // 2.0
    wire [14:0] v2073; shift_adder #(13, 13, 1, 1, 15, 2, 0) op_2073 (v645[12:0], v673[12:0], v2073[14:0]); // 2.0
    wire [19:0] v2074; shift_adder #(18, 19, 1, 1, 20, 1, 0) op_2074 (v286[17:0], v376[18:0], v2074[19:0]); // 2.0
    wire [13:0] v2075; shift_adder #(11, 11, 1, 1, 14, 3, 1) op_2075 (v140[10:0], v289[10:0], v2075[13:0]); // 2.0
    wire [13:0] v2076; shift_adder #(12, 11, 1, 1, 14, 3, 0) op_2076 (v397[11:0], v171[10:0], v2076[13:0]); // 2.0
    wire [11:0] v2077; shift_adder #(11, 10, 1, 1, 12, -1, 1) op_2077 (v208[10:0], v428[9:0], v2077[11:0]); // 2.0
    wire [12:0] v2078; shift_adder #(12, 12, 1, 1, 13, 1, 0) op_2078 (v239[11:0], v347[11:0], v2078[12:0]); // 2.0
    wire [14:0] v2079; shift_adder #(11, 15, 1, 1, 15, -1, 0) op_2079 (v269[10:0], v674[14:0], v2079[14:0]); // 2.0
    wire [15:0] v2080; shift_adder #(15, 11, 1, 1, 16, 4, 0) op_2080 (v649[14:0], v182[10:0], v2080[15:0]); // 2.0
    wire [12:0] v2081; shift_adder #(11, 12, 1, 1, 13, -2, 0) op_2081 (v675[10:0], v239[11:0], v2081[12:0]); // 2.0
    wire [13:0] v2082; shift_adder #(11, 13, 1, 1, 14, -2, 0) op_2082 (v676[10:0], v326[12:0], v2082[13:0]); // 2.0
    wire [11:0] v2083; shift_adder #(11, 11, 1, 1, 12, 0, 0) op_2083 (v284[10:0], v671[10:0], v2083[11:0]); // 2.0
    wire [12:0] v2084; shift_adder #(10, 11, 1, 1, 13, -3, 0) op_2084 (v263[9:0], v367[10:0], v2084[12:0]); // 2.0
    wire [11:0] v2085; shift_adder #(11, 10, 1, 1, 12, 1, 0) op_2085 (v165[10:0], v466[9:0], v2085[11:0]); // 2.0
    wire [11:0] v2086; shift_adder #(11, 11, 1, 1, 12, -1, 0) op_2086 (v497[10:0], v270[10:0], v2086[11:0]); // 2.0
    wire [30:0] v2087; shift_adder #(8, 10, 1, 1, 31, 21, 0) op_2087 (v65[7:0], v542[9:0], v2087[30:0]); // 2.0
    wire [15:0] v2088; shift_adder #(10, 16, 1, 1, 16, -2, 0) op_2088 (v260[9:0], v504[15:0], v2088[15:0]); // 2.0
    wire [21:0] v2089; shift_adder #(11, 21, 1, 1, 22, -10, 0) op_2089 (v324[10:0], v599[20:0], v2089[21:0]); // 2.0
    wire [12:0] v2090; shift_adder #(9, 9, 1, 1, 13, -3, 1) op_2090 (v401[8:0], v401[8:0], v2090[12:0]); // 2.0
    wire [13:0] v2091; shift_adder #(11, 12, 1, 1, 14, 2, 1) op_2091 (v277[10:0], v288[11:0], v2091[13:0]); // 2.0
    wire [34:0] v2092; shift_adder #(11, 10, 1, 1, 35, 25, 1) op_2092 (v275[10:0], v643[9:0], v2092[34:0]); // 2.0
    wire [16:0] v2093; shift_adder #(14, 17, 1, 1, 17, -2, 0) op_2093 (v410[13:0], v677[16:0], v2093[16:0]); // 2.0
    wire [11:0] v2094; shift_adder #(10, 11, 1, 1, 12, -1, 0) op_2094 (v678[9:0], v679[10:0], v2094[11:0]); // 2.0
    wire [10:0] v2095; shift_adder #(8, 11, 1, 1, 11, -1, 0) op_2095 (v73[7:0], v334[10:0], v2095[10:0]); // 2.0
    wire [23:0] v2096; shift_adder #(8, 24, 1, 1, 24, -1, 1) op_2096 (v125[7:0], v680[23:0], v2096[23:0]); // 2.0
    wire [27:0] v2097; shift_adder #(28, 18, 1, 1, 28, 8, 0) op_2097 (v618[27:0], v681[17:0], v2097[27:0]); // 2.0
    wire [12:0] v2098; shift_adder #(12, 10, 1, 1, 13, -1, 1) op_2098 (v357[11:0], v548[9:0], v2098[12:0]); // 2.0
    wire [14:0] v2099; shift_adder #(12, 12, 1, 1, 15, -3, 1) op_2099 (v438[11:0], v438[11:0], v2099[14:0]); // 2.0
    wire [12:0] v2100; shift_adder #(11, 12, 1, 1, 13, 1, 0) op_2100 (v298[10:0], v227[11:0], v2100[12:0]); // 2.0
    wire [13:0] v2101; shift_adder #(11, 12, 1, 1, 14, -3, 0) op_2101 (v671[10:0], v204[11:0], v2101[13:0]); // 2.0
    wire [10:0] v2102; shift_adder #(11, 9, 1, 1, 11, 0, 0) op_2102 (v176[10:0], v477[8:0], v2102[10:0]); // 2.0
    wire [25:0] v2103; shift_adder #(11, 11, 1, 1, 26, 15, 1) op_2103 (v141[10:0], v201[10:0], v2103[25:0]); // 2.0
    wire [9:0] v2104; shift_adder #(8, 9, 1, 1, 10, 0, 0) op_2104 (v107[7:0], v368[8:0], v2104[9:0]); // 2.0
    wire [14:0] v2105; shift_adder #(11, 12, 1, 1, 15, 3, 1) op_2105 (v287[10:0], v339[11:0], v2105[14:0]); // 2.0
    wire [14:0] v2106; shift_adder #(11, 12, 1, 1, 15, -4, 0) op_2106 (v162[10:0], v247[11:0], v2106[14:0]); // 2.0
    wire [11:0] v2107; shift_adder #(11, 9, 1, 1, 12, -1, 0) op_2107 (v176[10:0], v230[8:0], v2107[11:0]); // 2.0
    wire [11:0] v2108; shift_adder #(11, 12, 1, 1, 12, 0, 0) op_2108 (v420[10:0], v387[11:0], v2108[11:0]); // 2.0
    wire [14:0] v2109; shift_adder #(15, 12, 1, 1, 15, 2, 0) op_2109 (v630[14:0], v214[11:0], v2109[14:0]); // 2.0
    wire [13:0] v2110; shift_adder #(8, 11, 1, 1, 14, -5, 0) op_2110 (v64[7:0], v659[10:0], v2110[13:0]); // 2.0
    wire [14:0] v2111; shift_adder #(11, 11, 1, 1, 15, 4, 0) op_2111 (v135[10:0], v201[10:0], v2111[14:0]); // 2.0
    wire [16:0] v2112; shift_adder #(8, 10, 1, 1, 17, -8, 1) op_2112 (v116[7:0], v549[9:0], v2112[16:0]); // 2.0
    wire [14:0] v2113; shift_adder #(10, 14, 1, 1, 15, 1, 0) op_2113 (v282[9:0], v394[13:0], v2113[14:0]); // 2.0
    wire [22:0] v2114; shift_adder #(8, 11, 1, 1, 23, -14, 1) op_2114 (v111[7:0], v154[10:0], v2114[22:0]); // 2.0
    wire [13:0] v2115; shift_adder #(12, 12, 1, 1, 14, 2, 0) op_2115 (v552[11:0], v614[11:0], v2115[13:0]); // 2.0
    wire [11:0] v2116; shift_adder #(11, 11, 1, 1, 12, 1, 0) op_2116 (v157[10:0], v150[10:0], v2116[11:0]); // 2.0
    wire [14:0] v2117; shift_adder #(11, 13, 1, 1, 15, -4, 0) op_2117 (v173[10:0], v192[12:0], v2117[14:0]); // 2.0
    wire [13:0] v2118; shift_adder #(11, 12, 1, 1, 14, 2, 1) op_2118 (v276[10:0], v382[11:0], v2118[13:0]); // 2.0
    wire [18:0] v2119; shift_adder #(11, 19, 1, 1, 19, -3, 0) op_2119 (v574[10:0], v547[18:0], v2119[18:0]); // 2.0
    wire [20:0] v2120; shift_adder #(20, 18, 1, 1, 21, 3, 0) op_2120 (v515[19:0], v535[17:0], v2120[20:0]); // 2.0
    wire [29:0] v2121; shift_adder #(11, 18, 1, 1, 30, 12, 0) op_2121 (v161[10:0], v682[17:0], v2121[29:0]); // 2.0
    wire [13:0] v2122; shift_adder #(11, 13, 1, 1, 14, -2, 0) op_2122 (v518[10:0], v344[12:0], v2122[13:0]); // 2.0
    wire [10:0] v2123; shift_adder #(8, 11, 1, 1, 11, 0, 1) op_2123 (v125[7:0], v353[10:0], v2123[10:0]); // 2.0
    wire [11:0] v2124; shift_adder #(8, 12, 1, 1, 12, -2, 0) op_2124 (v64[7:0], v146[11:0], v2124[11:0]); // 2.0
    wire [34:0] v2125; shift_adder #(12, 35, 1, 1, 35, -22, 0) op_2125 (v438[11:0], v683[34:0], v2125[34:0]); // 2.0
    wire [12:0] v2126; shift_adder #(10, 12, 1, 1, 13, -2, 0) op_2126 (v470[9:0], v389[11:0], v2126[12:0]); // 2.0
    wire [12:0] v2127; shift_adder #(10, 11, 1, 1, 13, -3, 0) op_2127 (v450[9:0], v215[10:0], v2127[12:0]); // 2.0
    wire [32:0] v2128; shift_adder #(11, 32, 1, 1, 33, -21, 0) op_2128 (v255[10:0], v684[31:0], v2128[32:0]); // 2.0
    wire [10:0] v2129; shift_adder #(10, 11, 1, 1, 11, 0, 0) op_2129 (v527[9:0], v685[10:0], v2129[10:0]); // 2.0
    wire [11:0] v2130; shift_adder #(12, 11, 1, 1, 12, 0, 0) op_2130 (v521[11:0], v232[10:0], v2130[11:0]); // 2.0
    wire [19:0] v2131; shift_adder #(13, 17, 1, 1, 20, -7, 0) op_2131 (v573[12:0], v335[16:0], v2131[19:0]); // 2.0
    wire [12:0] v2132; shift_adder #(12, 11, 1, 1, 13, 1, 0) op_2132 (v462[11:0], v218[10:0], v2132[12:0]); // 2.0
    wire [12:0] v2133; shift_adder #(12, 12, 1, 1, 13, 0, 0) op_2133 (v686[11:0], v363[11:0], v2133[12:0]); // 2.0
    wire [13:0] v2134; shift_adder #(11, 11, 1, 1, 14, -3, 1) op_2134 (v177[10:0], v361[10:0], v2134[13:0]); // 2.0
    wire [11:0] v2135; shift_adder #(11, 11, 1, 1, 12, 1, 0) op_2135 (v175[10:0], v319[10:0], v2135[11:0]); // 2.0
    wire [13:0] v2136; shift_adder #(13, 13, 1, 1, 14, -1, 0) op_2136 (v578[12:0], v598[12:0], v2136[13:0]); // 2.0
    wire [11:0] v2137; shift_adder #(11, 11, 1, 1, 12, 0, 0) op_2137 (v303[10:0], v228[10:0], v2137[11:0]); // 2.0
    wire [25:0] v2138; shift_adder #(24, 9, 1, 1, 26, 16, 0) op_2138 (v680[23:0], v568[8:0], v2138[25:0]); // 2.0
    wire [12:0] v2139; shift_adder #(12, 11, 1, 1, 13, -1, 0) op_2139 (v321[11:0], v284[10:0], v2139[12:0]); // 2.0
    wire [17:0] v2140; shift_adder #(11, 11, 1, 1, 18, -7, 0) op_2140 (v229[10:0], v270[10:0], v2140[17:0]); // 2.0
    wire [12:0] v2141; shift_adder #(8, 12, 1, 1, 13, 1, 0) op_2141 (v79[7:0], v398[11:0], v2141[12:0]); // 2.0
    wire [17:0] v2142; shift_adder #(14, 16, 1, 1, 18, -4, 0) op_2142 (v687[13:0], v240[15:0], v2142[17:0]); // 2.0
    wire [13:0] v2143; shift_adder #(8, 12, 1, 1, 14, -5, 0) op_2143 (v80[7:0], v434[11:0], v2143[13:0]); // 2.0
    wire [21:0] v2144; shift_adder #(22, 18, 1, 1, 22, 2, 0) op_2144 (v656[21:0], v286[17:0], v2144[21:0]); // 2.0
    wire [17:0] v2145; shift_adder #(11, 11, 1, 1, 18, -7, 0) op_2145 (v212[10:0], v430[10:0], v2145[17:0]); // 2.0
    wire [13:0] v2146; shift_adder #(9, 11, 1, 1, 14, -4, 0) op_2146 (v441[8:0], v206[10:0], v2146[13:0]); // 2.0
    wire [13:0] v2147; shift_adder #(11, 12, 1, 1, 14, -3, 0) op_2147 (v518[10:0], v257[11:0], v2147[13:0]); // 2.0
    wire [29:0] v2148; shift_adder #(11, 23, 1, 1, 30, -19, 0) op_2148 (v211[10:0], v580[22:0], v2148[29:0]); // 2.0
    wire [20:0] v2149; shift_adder #(13, 21, 1, 1, 21, -7, 0) op_2149 (v198[12:0], v364[20:0], v2149[20:0]); // 2.0
    wire [15:0] v2150; shift_adder #(11, 11, 1, 1, 16, -5, 1) op_2150 (v188[10:0], v212[10:0], v2150[15:0]); // 2.0
    wire [23:0] v2151; shift_adder #(8, 12, 1, 1, 24, 12, 0) op_2151 (v95[7:0], v550[11:0], v2151[23:0]); // 2.0
    wire [11:0] v2152; shift_adder #(9, 11, 1, 1, 12, -1, 0) op_2152 (v637[8:0], v165[10:0], v2152[11:0]); // 2.0
    wire [28:0] v2153; shift_adder #(11, 12, 1, 1, 29, -18, 1) op_2153 (v133[10:0], v280[11:0], v2153[28:0]); // 2.0
    wire [11:0] v2154; shift_adder #(9, 11, 1, 1, 12, 1, 0) op_2154 (v663[8:0], v688[10:0], v2154[11:0]); // 2.0
    wire [16:0] v2155; shift_adder #(13, 13, 1, 1, 17, 4, 0) op_2155 (v272[12:0], v476[12:0], v2155[16:0]); // 2.0
    wire [12:0] v2156; shift_adder #(12, 11, 1, 1, 13, 2, 0) op_2156 (v339[11:0], v255[10:0], v2156[12:0]); // 2.0
    wire [16:0] v2157; shift_adder #(11, 17, 1, 1, 17, -4, 0) op_2157 (v241[10:0], v689[16:0], v2157[16:0]); // 2.0
    wire [11:0] v2158; shift_adder #(11, 11, 1, 1, 12, 0, 0) op_2158 (v425[10:0], v269[10:0], v2158[11:0]); // 2.0
    wire [14:0] v2159; shift_adder #(11, 13, 1, 1, 15, -4, 0) op_2159 (v338[10:0], v534[12:0], v2159[14:0]); // 2.0
    wire [15:0] v2160; shift_adder #(15, 11, 1, 1, 16, 5, 0) op_2160 (v690[14:0], v228[10:0], v2160[15:0]); // 2.0
    wire [18:0] v2161; shift_adder #(11, 19, 1, 1, 19, -6, 0) op_2161 (v219[10:0], v640[18:0], v2161[18:0]); // 2.0
    wire [11:0] v2162; shift_adder #(11, 12, 1, 1, 12, 0, 0) op_2162 (v328[10:0], v691[11:0], v2162[11:0]); // 2.0
    wire [33:0] v2163; shift_adder #(11, 10, 1, 1, 34, -23, 1) op_2163 (v136[10:0], v366[9:0], v2163[33:0]); // 2.0
    wire [10:0] v2164; shift_adder #(11, 10, 1, 1, 11, 0, 0) op_2164 (v692[10:0], v252[9:0], v2164[10:0]); // 2.0
    wire [11:0] v2165; shift_adder #(11, 11, 1, 1, 12, 1, 0) op_2165 (v505[10:0], v430[10:0], v2165[11:0]); // 2.0
    wire [34:0] v2166; shift_adder #(9, 8, 1, 1, 35, 26, 1) op_2166 (v256[8:0], v84[7:0], v2166[34:0]); // 2.0
    wire [12:0] v2167; shift_adder #(12, 9, 1, 1, 13, 3, 0) op_2167 (v357[11:0], v693[8:0], v2167[12:0]); // 2.0
    wire [11:0] v2168; shift_adder #(11, 11, 1, 1, 12, -1, 0) op_2168 (v251[10:0], v163[10:0], v2168[11:0]); // 2.0
    wire [16:0] v2169; shift_adder #(17, 11, 1, 1, 17, 4, 0) op_2169 (v551[16:0], v141[10:0], v2169[16:0]); // 2.0
    wire [12:0] v2170; shift_adder #(11, 11, 1, 1, 13, 2, 0) op_2170 (v134[10:0], v197[10:0], v2170[12:0]); // 2.0
    wire [12:0] v2171; shift_adder #(12, 12, 1, 1, 13, -1, 1) op_2171 (v521[11:0], v579[11:0], v2171[12:0]); // 2.0
    wire [19:0] v2172; shift_adder #(11, 11, 1, 1, 20, 9, 1) op_2172 (v270[10:0], v497[10:0], v2172[19:0]); // 2.0
    wire [16:0] v2173; shift_adder #(11, 12, 1, 1, 17, -6, 1) op_2173 (v283[10:0], v321[11:0], v2173[16:0]); // 2.0
    wire [12:0] v2174; shift_adder #(11, 11, 1, 1, 13, -2, 0) op_2174 (v694[10:0], v413[10:0], v2174[12:0]); // 2.0
    wire [14:0] v2175; shift_adder #(11, 15, 1, 1, 15, -3, 0) op_2175 (v181[10:0], v695[14:0], v2175[14:0]); // 2.0
    wire [12:0] v2176; shift_adder #(9, 11, 1, 1, 13, -3, 0) op_2176 (v637[8:0], v696[10:0], v2176[12:0]); // 2.0
    wire [12:0] v2177; shift_adder #(13, 10, 1, 1, 13, 1, 0) op_2177 (v506[12:0], v468[9:0], v2177[12:0]); // 2.0
    wire [13:0] v2178; shift_adder #(13, 11, 1, 1, 14, 2, 0) op_2178 (v451[12:0], v195[10:0], v2178[13:0]); // 2.0
    wire [11:0] v2179; shift_adder #(10, 12, 1, 1, 12, -1, 0) op_2179 (v468[9:0], v265[11:0], v2179[11:0]); // 2.0
    wire [11:0] v2180; shift_adder #(10, 12, 1, 1, 12, 0, 0) op_2180 (v565[9:0], v502[11:0], v2180[11:0]); // 2.0
    wire [23:0] v2181; shift_adder #(8, 12, 1, 1, 24, 12, 0) op_2181 (v74[7:0], v174[11:0], v2181[23:0]); // 2.0
    wire [17:0] v2182; shift_adder #(17, 11, 1, 1, 18, 7, 0) op_2182 (v348[16:0], v228[10:0], v2182[17:0]); // 2.0
    wire [9:0] v2183; shift_adder #(8, 9, 1, 1, 10, -1, 1) op_2183 (v103[7:0], v360[8:0], v2183[9:0]); // 2.0
    wire [12:0] v2184; shift_adder #(11, 11, 1, 1, 13, 2, 0) op_2184 (v245[10:0], v212[10:0], v2184[12:0]); // 2.0
    wire [15:0] v2185; shift_adder #(8, 11, 1, 1, 16, -7, 1) op_2185 (v121[7:0], v234[10:0], v2185[15:0]); // 2.0
    wire [13:0] v2186; shift_adder #(8, 11, 1, 1, 14, -5, 0) op_2186 (v105[7:0], v250[10:0], v2186[13:0]); // 2.0
    wire [16:0] v2187; shift_adder #(15, 11, 1, 1, 17, 6, 0) op_2187 (v697[14:0], v181[10:0], v2187[16:0]); // 2.0
    wire [11:0] v2188; shift_adder #(11, 11, 1, 1, 12, 0, 0) op_2188 (v168[10:0], v299[10:0], v2188[11:0]); // 2.0
    wire [14:0] v2189; shift_adder #(11, 10, 1, 1, 15, 5, 1) op_2189 (v157[10:0], v291[9:0], v2189[14:0]); // 2.0
    wire [11:0] v2190; shift_adder #(11, 12, 1, 1, 12, 0, 0) op_2190 (v671[10:0], v325[11:0], v2190[11:0]); // 2.0
    wire [35:0] v2191; shift_adder #(14, 8, 1, 1, 36, 27, 1) op_2191 (v698[13:0], v126[7:0], v2191[35:0]); // 2.0
    wire [12:0] v2192; shift_adder #(12, 9, 1, 1, 13, 3, 0) op_2192 (v582[11:0], v302[8:0], v2192[12:0]); // 2.0
    wire [18:0] v2193; shift_adder #(9, 18, 1, 1, 19, -8, 0) op_2193 (v138[8:0], v494[17:0], v2193[18:0]); // 2.0
    wire [10:0] v2194; shift_adder #(8, 10, 1, 1, 11, -1, 0) op_2194 (v101[7:0], v592[9:0], v2194[10:0]); // 2.0
    wire [10:0] v2195; shift_adder #(10, 11, 1, 1, 11, 0, 0) op_2195 (v699[9:0], v168[10:0], v2195[10:0]); // 2.0
    wire [12:0] v2196; shift_adder #(13, 11, 1, 1, 13, 1, 0) op_2196 (v645[12:0], v173[10:0], v2196[12:0]); // 2.0
    wire [18:0] v2197; shift_adder #(8, 11, 1, 1, 19, -10, 1) op_2197 (v95[7:0], v216[10:0], v2197[18:0]); // 2.0
    wire [16:0] v2198; shift_adder #(15, 10, 1, 1, 17, 6, 0) op_2198 (v700[14:0], v273[9:0], v2198[16:0]); // 2.0
    wire [13:0] v2199; shift_adder #(11, 11, 1, 1, 14, 3, 1) op_2199 (v301[10:0], v246[10:0], v2199[13:0]); // 2.0
    wire [11:0] v2200; shift_adder #(12, 9, 1, 1, 12, 1, 0) op_2200 (v552[11:0], v230[8:0], v2200[11:0]); // 2.0
    wire [14:0] v2201; shift_adder #(11, 13, 1, 1, 15, -4, 0) op_2201 (v140[10:0], v598[12:0], v2201[14:0]); // 2.0
    wire [10:0] v2202; shift_adder #(10, 10, 1, 1, 11, 0, 0) op_2202 (v435[9:0], v254[9:0], v2202[10:0]); // 2.0
    wire [25:0] v2203; shift_adder #(11, 12, 1, 1, 26, 14, 1) op_2203 (v154[10:0], v180[11:0], v2203[25:0]); // 2.0
    wire [20:0] v2204; shift_adder #(11, 11, 1, 1, 21, -10, 0) op_2204 (v284[10:0], v197[10:0], v2204[20:0]); // 2.0
    wire [13:0] v2205; shift_adder #(12, 13, 1, 1, 14, -1, 0) op_2205 (v540[11:0], v198[12:0], v2205[13:0]); // 2.0
    wire [20:0] v2206; shift_adder #(11, 14, 1, 1, 21, -10, 1) op_2206 (v375[10:0], v571[13:0], v2206[20:0]); // 2.0
    wire [13:0] v2207; shift_adder #(13, 11, 1, 1, 14, 2, 0) op_2207 (v416[12:0], v701[10:0], v2207[13:0]); // 2.0
    wire [17:0] v2208; shift_adder #(11, 12, 1, 1, 18, 6, 0) op_2208 (v393[10:0], v202[11:0], v2208[17:0]); // 2.0
    wire [15:0] v2209; shift_adder #(11, 12, 1, 1, 16, 4, 0) op_2209 (v379[10:0], v462[11:0], v2209[15:0]); // 2.0
    wire [13:0] v2210; shift_adder #(11, 11, 1, 1, 14, -3, 0) op_2210 (v702[10:0], v345[10:0], v2210[13:0]); // 2.0
    wire [15:0] v2211; shift_adder #(12, 15, 1, 1, 16, -3, 0) op_2211 (v380[11:0], v703[14:0], v2211[15:0]); // 2.0
    wire [20:0] v2212; shift_adder #(21, 11, 1, 1, 21, 9, 0) op_2212 (v364[20:0], v320[10:0], v2212[20:0]); // 2.0
    wire [11:0] v2213; shift_adder #(11, 11, 1, 1, 12, 0, 0) op_2213 (v144[10:0], v418[10:0], v2213[11:0]); // 2.0
    wire [12:0] v2214; shift_adder #(12, 11, 1, 1, 13, 2, 0) op_2214 (v392[11:0], v140[10:0], v2214[12:0]); // 2.0
    wire [12:0] v2215; shift_adder #(8, 12, 1, 1, 13, 1, 0) op_2215 (v126[7:0], v184[11:0], v2215[12:0]); // 2.0
    wire [17:0] v2216; shift_adder #(10, 17, 1, 1, 18, -7, 0) op_2216 (v291[9:0], v689[16:0], v2216[17:0]); // 2.0
    wire [13:0] v2217; shift_adder #(12, 10, 1, 1, 14, 3, 0) op_2217 (v257[11:0], v468[9:0], v2217[13:0]); // 2.0
    wire [12:0] v2218; shift_adder #(13, 10, 1, 1, 13, 0, 1) op_2218 (v601[12:0], v584[9:0], v2218[12:0]); // 2.0
    wire [11:0] v2219; shift_adder #(10, 11, 1, 1, 12, 1, 0) op_2219 (v704[9:0], v287[10:0], v2219[11:0]); // 2.0
    wire [24:0] v2220; shift_adder #(11, 25, 1, 1, 25, -9, 0) op_2220 (v266[10:0], v595[24:0], v2220[24:0]); // 2.0
    wire [14:0] v2221; shift_adder #(12, 15, 1, 1, 15, -2, 0) op_2221 (v521[11:0], v465[14:0], v2221[14:0]); // 2.0
    wire [13:0] v2222; shift_adder #(11, 11, 1, 1, 14, -3, 0) op_2222 (v688[10:0], v200[10:0], v2222[13:0]); // 2.0
    wire [13:0] v2223; shift_adder #(12, 12, 1, 1, 14, 2, 0) op_2223 (v447[11:0], v357[11:0], v2223[13:0]); // 2.0
    wire [16:0] v2224; shift_adder #(13, 17, 1, 1, 17, -2, 1) op_2224 (v654[12:0], v348[16:0], v2224[16:0]); // 2.0
    wire [12:0] v2225; shift_adder #(11, 11, 1, 1, 13, -2, 0) op_2225 (v283[10:0], v172[10:0], v2225[12:0]); // 2.0
    wire [16:0] v2226; shift_adder #(11, 11, 1, 1, 17, 6, 0) op_2226 (v211[10:0], v162[10:0], v2226[16:0]); // 2.0
    wire [11:0] v2227; shift_adder #(10, 11, 1, 1, 12, 1, 0) op_2227 (v705[9:0], v352[10:0], v2227[11:0]); // 2.0
    wire [29:0] v2228; shift_adder #(10, 8, 1, 1, 30, 21, 1) op_2228 (v273[9:0], v125[7:0], v2228[29:0]); // 2.0
    wire [11:0] v2229; shift_adder #(11, 11, 1, 1, 12, -1, 0) op_2229 (v358[10:0], v233[10:0], v2229[11:0]); // 2.0
    wire [17:0] v2230; shift_adder #(8, 11, 1, 1, 18, -9, 0) op_2230 (v99[7:0], v141[10:0], v2230[17:0]); // 2.0
    wire [11:0] v2231; shift_adder #(11, 11, 1, 1, 12, 1, 0) op_2231 (v294[10:0], v218[10:0], v2231[11:0]); // 2.0
    wire [14:0] v2232; shift_adder #(15, 13, 1, 1, 15, 0, 0) op_2232 (v706[14:0], v534[12:0], v2232[14:0]); // 2.0
    wire [11:0] v2233; shift_adder #(9, 10, 1, 1, 12, 2, 0) op_2233 (v503[8:0], v707[9:0], v2233[11:0]); // 2.0
    wire [10:0] v2234; shift_adder #(8, 10, 1, 1, 11, -1, 0) op_2234 (v75[7:0], v366[9:0], v2234[10:0]); // 2.0
    wire [12:0] v2235; shift_adder #(11, 11, 1, 1, 13, 2, 0) op_2235 (v218[10:0], v245[10:0], v2235[12:0]); // 2.0
    wire [12:0] v2236; shift_adder #(12, 9, 1, 1, 13, 2, 0) op_2236 (v292[11:0], v322[8:0], v2236[12:0]); // 2.0
    wire [14:0] v2237; shift_adder #(13, 13, 1, 1, 15, 2, 0) op_2237 (v346[12:0], v492[12:0], v2237[14:0]); // 2.0
    wire [11:0] v2238; shift_adder #(8, 11, 1, 1, 12, -3, 1) op_2238 (v79[7:0], v200[10:0], v2238[11:0]); // 2.0
    wire [33:0] v2239; shift_adder #(17, 10, 1, 1, 34, -17, 1) op_2239 (v551[16:0], v260[9:0], v2239[33:0]); // 2.0
    wire [12:0] v2240; shift_adder #(12, 11, 1, 1, 13, 1, 0) op_2240 (v579[11:0], v478[10:0], v2240[12:0]); // 2.0
    wire [10:0] v2241; shift_adder #(11, 9, 1, 1, 11, 0, 0) op_2241 (v708[10:0], v302[8:0], v2241[10:0]); // 2.0
    wire [13:0] v2242; shift_adder #(13, 11, 1, 1, 14, 2, 0) op_2242 (v449[12:0], v211[10:0], v2242[13:0]); // 2.0
    wire [14:0] v2243; shift_adder #(11, 12, 1, 1, 15, -4, 1) op_2243 (v162[10:0], v224[11:0], v2243[14:0]); // 2.0
    wire [13:0] v2244; shift_adder #(14, 12, 1, 1, 14, 1, 0) op_2244 (v514[13:0], v709[11:0], v2244[13:0]); // 2.0
    wire [11:0] v2245; shift_adder #(11, 10, 1, 1, 12, -1, 0) op_2245 (v300[10:0], v459[9:0], v2245[11:0]); // 2.0
    wire [15:0] v2246; shift_adder #(9, 15, 1, 1, 16, -6, 0) op_2246 (v486[8:0], v313[14:0], v2246[15:0]); // 2.0
    wire [11:0] v2247; shift_adder #(11, 9, 1, 1, 12, 2, 0) op_2247 (v153[10:0], v256[8:0], v2247[11:0]); // 2.0
    wire [17:0] v2248; shift_adder #(11, 16, 1, 1, 18, -7, 0) op_2248 (v140[10:0], v710[15:0], v2248[17:0]); // 2.0
    wire [17:0] v2249; shift_adder #(10, 12, 1, 1, 18, -8, 0) op_2249 (v584[9:0], v357[11:0], v2249[17:0]); // 2.0
    wire [11:0] v2250; shift_adder #(11, 9, 1, 1, 12, -1, 0) op_2250 (v211[10:0], v503[8:0], v2250[11:0]); // 2.0
    wire [11:0] v2251; shift_adder #(11, 11, 1, 1, 12, -1, 0) op_2251 (v659[10:0], v147[10:0], v2251[11:0]); // 2.0
    wire [11:0] v2252; shift_adder #(11, 11, 1, 1, 12, 1, 0) op_2252 (v341[10:0], v300[10:0], v2252[11:0]); // 2.0
    wire [15:0] v2253; shift_adder #(14, 16, 1, 1, 16, -1, 0) op_2253 (v342[13:0], v711[15:0], v2253[15:0]); // 2.0
    wire [11:0] v2254; shift_adder #(10, 11, 1, 1, 12, -1, 0) op_2254 (v170[9:0], v134[10:0], v2254[11:0]); // 2.0
    wire [19:0] v2255; shift_adder #(11, 11, 1, 1, 20, 9, 1) op_2255 (v223[10:0], v206[10:0], v2255[19:0]); // 2.0
    wire [11:0] v2256; shift_adder #(11, 12, 1, 1, 12, 0, 0) op_2256 (v199[10:0], v540[11:0], v2256[11:0]); // 2.0
    wire [25:0] v2257; shift_adder #(15, 26, 1, 1, 26, -9, 0) op_2257 (v465[14:0], v525[25:0], v2257[25:0]); // 2.0
    wire [12:0] v2258; shift_adder #(8, 11, 1, 1, 13, -4, 1) op_2258 (v120[7:0], v155[10:0], v2258[12:0]); // 2.0
    wire [12:0] v2259; shift_adder #(9, 11, 1, 1, 13, -3, 0) op_2259 (v568[8:0], v179[10:0], v2259[12:0]); // 2.0
    wire [10:0] v2260; shift_adder #(9, 10, 1, 1, 11, -1, 1) op_2260 (v302[8:0], v282[9:0], v2260[10:0]); // 2.0
    wire [23:0] v2261; shift_adder #(11, 11, 1, 1, 24, -13, 1) op_2261 (v396[10:0], v268[10:0], v2261[23:0]); // 2.0
    wire [38:0] v2262; shift_adder #(11, 12, 1, 1, 39, -28, 1) op_2262 (v134[10:0], v541[11:0], v2262[38:0]); // 2.0
    wire [35:0] v2263; shift_adder #(10, 8, 1, 1, 36, 27, 1) op_2263 (v705[9:0], v77[7:0], v2263[35:0]); // 2.0
    wire [12:0] v2264; shift_adder #(11, 11, 1, 1, 13, -2, 0) op_2264 (v188[10:0], v276[10:0], v2264[12:0]); // 2.0
    wire [13:0] v2265; shift_adder #(11, 11, 1, 1, 14, 3, 0) op_2265 (v317[10:0], v319[10:0], v2265[13:0]); // 2.0
    wire [15:0] v2266; shift_adder #(11, 12, 1, 1, 16, -5, 0) op_2266 (v712[10:0], v553[11:0], v2266[15:0]); // 2.0
    wire [14:0] v2267; shift_adder #(11, 11, 1, 1, 15, -4, 0) op_2267 (v283[10:0], v233[10:0], v2267[14:0]); // 2.0
    wire [12:0] v2268; shift_adder #(8, 11, 1, 1, 13, -4, 0) op_2268 (v123[7:0], v203[10:0], v2268[12:0]); // 2.0
    wire [15:0] v2269; shift_adder #(13, 16, 1, 1, 16, -2, 0) op_2269 (v416[12:0], v504[15:0], v2269[15:0]); // 2.0
    wire [15:0] v2270; shift_adder #(15, 12, 1, 1, 16, 3, 0) op_2270 (v471[14:0], v365[11:0], v2270[15:0]); // 2.0
    wire [15:0] v2271; shift_adder #(8, 14, 1, 1, 16, -7, 1) op_2271 (v71[7:0], v483[13:0], v2271[15:0]); // 2.0
    wire [29:0] v2272; shift_adder #(11, 29, 1, 1, 30, -18, 0) op_2272 (v203[10:0], v713[28:0], v2272[29:0]); // 2.0
    wire [13:0] v2273; shift_adder #(11, 12, 1, 1, 14, -3, 1) op_2273 (v386[10:0], v541[11:0], v2273[13:0]); // 2.0
    wire [11:0] v2274; shift_adder #(11, 11, 1, 1, 12, 0, 0) op_2274 (v714[10:0], v574[10:0], v2274[11:0]); // 2.0
    wire [13:0] v2275; shift_adder #(13, 11, 1, 1, 14, 2, 0) op_2275 (v715[12:0], v268[10:0], v2275[13:0]); // 2.0
    wire [13:0] v2276; shift_adder #(10, 11, 1, 1, 14, -4, 0) op_2276 (v716[9:0], v242[10:0], v2276[13:0]); // 2.0
    wire [16:0] v2277; shift_adder #(11, 11, 1, 1, 17, 6, 1) op_2277 (v172[10:0], v334[10:0], v2277[16:0]); // 2.0
    wire [26:0] v2278; shift_adder #(11, 12, 1, 1, 27, 15, 0) op_2278 (v178[10:0], v614[11:0], v2278[26:0]); // 2.0
    wire [20:0] v2279; shift_adder #(11, 9, 1, 1, 21, 12, 0) op_2279 (v420[10:0], v369[8:0], v2279[20:0]); // 2.0
    wire [16:0] v2280; shift_adder #(17, 10, 1, 1, 17, 4, 0) op_2280 (v615[16:0], v717[9:0], v2280[16:0]); // 2.0
    wire [12:0] v2281; shift_adder #(11, 11, 1, 1, 13, -2, 0) op_2281 (v353[10:0], v275[10:0], v2281[12:0]); // 2.0
    wire [13:0] v2282; shift_adder #(13, 9, 1, 1, 14, 4, 0) op_2282 (v718[12:0], v309[8:0], v2282[13:0]); // 2.0
    wire [11:0] v2283; shift_adder #(11, 11, 1, 1, 12, -1, 0) op_2283 (v154[10:0], v234[10:0], v2283[11:0]); // 2.0
    wire [12:0] v2284; shift_adder #(11, 11, 1, 1, 13, -2, 0) op_2284 (v250[10:0], v714[10:0], v2284[12:0]); // 2.0
    wire [12:0] v2285; shift_adder #(11, 12, 1, 1, 13, 1, 0) op_2285 (v144[10:0], v719[11:0], v2285[12:0]); // 2.0
    wire [11:0] v2286; shift_adder #(11, 12, 1, 1, 12, 0, 1) op_2286 (v299[10:0], v387[11:0], v2286[11:0]); // 2.0
    wire [13:0] v2287; shift_adder #(10, 9, 1, 1, 14, 4, 0) op_2287 (v510[9:0], v302[8:0], v2287[13:0]); // 2.0
    wire [13:0] v2288; shift_adder #(12, 13, 1, 1, 14, -1, 0) op_2288 (v347[11:0], v416[12:0], v2288[13:0]); // 2.0
    wire [17:0] v2289; shift_adder #(11, 11, 1, 1, 18, 7, 0) op_2289 (v158[10:0], v213[10:0], v2289[17:0]); // 2.0
    wire [9:0] v2290; shift_adder #(8, 10, 1, 1, 10, 0, 0) op_2290 (v126[7:0], v610[9:0], v2290[9:0]); // 2.0
    wire [31:0] v2291; shift_adder #(8, 14, 1, 1, 32, 18, 1) op_2291 (v107[7:0], v290[13:0], v2291[31:0]); // 2.0
    wire [11:0] v2292; shift_adder #(11, 11, 1, 1, 12, 1, 0) op_2292 (v176[10:0], v215[10:0], v2292[11:0]); // 2.0
    wire [10:0] v2293; shift_adder #(8, 9, 1, 1, 11, -2, 1) op_2293 (v101[7:0], v221[8:0], v2293[10:0]); // 2.0
    wire [11:0] v2294; shift_adder #(11, 9, 1, 1, 12, 1, 0) op_2294 (v173[10:0], v621[8:0], v2294[11:0]); // 2.0
    wire [12:0] v2295; shift_adder #(12, 11, 1, 1, 13, 2, 0) op_2295 (v452[11:0], v259[10:0], v2295[12:0]); // 2.0
    wire [20:0] v2296; shift_adder #(11, 11, 1, 1, 21, -10, 0) op_2296 (v175[10:0], v175[10:0], v2296[20:0]); // 2.0
    wire [16:0] v2297; shift_adder #(12, 12, 1, 1, 17, 5, 0) op_2297 (v423[11:0], v288[11:0], v2297[16:0]); // 2.0
    wire [12:0] v2298; shift_adder #(11, 11, 1, 1, 13, -2, 1) op_2298 (v193[10:0], v150[10:0], v2298[12:0]); // 2.0
    wire [17:0] v2299; shift_adder #(18, 11, 1, 1, 18, 4, 0) op_2299 (v682[17:0], v317[10:0], v2299[17:0]); // 2.0
    wire [26:0] v2300; shift_adder #(27, 11, 1, 1, 27, 13, 0) op_2300 (v720[26:0], v246[10:0], v2300[26:0]); // 2.0
    wire [16:0] v2301; shift_adder #(16, 9, 1, 1, 17, 7, 0) op_2301 (v240[15:0], v556[8:0], v2301[16:0]); // 2.0
    wire [11:0] v2302; shift_adder #(11, 11, 1, 1, 12, 1, 0) op_2302 (v129[10:0], v721[10:0], v2302[11:0]); // 2.0
    wire [11:0] v2303; shift_adder #(10, 11, 1, 1, 12, -1, 0) op_2303 (v716[9:0], v139[10:0], v2303[11:0]); // 2.0
    wire [13:0] v2304; shift_adder #(11, 12, 1, 1, 14, -3, 0) op_2304 (v443[10:0], v382[11:0], v2304[13:0]); // 2.0
    wire [11:0] v2305; shift_adder #(11, 9, 1, 1, 12, 1, 0) op_2305 (v723[10:0], v620[8:0], v2305[11:0]); // 2.0
    wire [12:0] v2306; shift_adder #(11, 9, 1, 1, 13, 3, 0) op_2306 (v320[10:0], v724[8:0], v2306[12:0]); // 2.0
    wire [34:0] v2307; shift_adder #(34, 10, 1, 1, 35, 25, 0) op_2307 (v399[33:0], v435[9:0], v2307[34:0]); // 2.0
    wire [33:0] v2308; shift_adder #(22, 11, 1, 1, 34, -12, 1) op_2308 (v656[21:0], v577[10:0], v2308[33:0]); // 2.0
    wire [13:0] v2309; shift_adder #(14, 9, 1, 1, 14, 2, 0) op_2309 (v488[13:0], v467[8:0], v2309[13:0]); // 2.0
    wire [12:0] v2310; shift_adder #(13, 11, 1, 1, 13, 1, 0) op_2310 (v534[12:0], v274[10:0], v2310[12:0]); // 2.0
    wire [27:0] v2311; shift_adder #(8, 11, 1, 1, 28, -19, 1) op_2311 (v80[7:0], v185[10:0], v2311[27:0]); // 2.0
    wire [25:0] v2312; shift_adder #(12, 24, 1, 1, 26, -14, 0) op_2312 (v357[11:0], v725[23:0], v2312[25:0]); // 2.0
    wire [11:0] v2313; shift_adder #(11, 11, 1, 1, 12, -1, 0) op_2313 (v303[10:0], v185[10:0], v2313[11:0]); // 2.0
    wire [23:0] v2314; shift_adder #(8, 11, 1, 1, 24, -15, 1) op_2314 (v89[7:0], v155[10:0], v2314[23:0]); // 2.0
    wire [11:0] v2315; shift_adder #(11, 10, 1, 1, 12, -1, 0) op_2315 (v317[10:0], v366[9:0], v2315[11:0]); // 2.0
    wire [13:0] v2316; shift_adder #(12, 11, 1, 1, 14, 3, 0) op_2316 (v407[11:0], v379[10:0], v2316[13:0]); // 2.0
    wire [18:0] v2317; shift_adder #(11, 12, 1, 1, 19, 7, 1) op_2317 (v353[10:0], v473[11:0], v2317[18:0]); // 2.0
    wire [13:0] v2318; shift_adder #(10, 12, 1, 1, 14, -3, 0) op_2318 (v554[9:0], v629[11:0], v2318[13:0]); // 2.0
    wire [17:0] v2319; shift_adder #(11, 18, 1, 1, 18, -4, 0) op_2319 (v155[10:0], v633[17:0], v2319[17:0]); // 2.0
    wire [15:0] v2320; shift_adder #(11, 11, 1, 1, 16, 5, 0) op_2320 (v232[10:0], v201[10:0], v2320[15:0]); // 2.0
    wire [10:0] v2321; shift_adder #(9, 10, 1, 1, 11, -1, 0) op_2321 (v384[8:0], v222[9:0], v2321[10:0]); // 2.0
    wire [18:0] v2322; shift_adder #(16, 19, 1, 1, 19, -2, 0) op_2322 (v240[15:0], v315[18:0], v2322[18:0]); // 2.0
    wire [14:0] v2323; shift_adder #(11, 12, 1, 1, 15, 3, 1) op_2323 (v374[10:0], v337[11:0], v2323[14:0]); // 2.0
    wire [17:0] v2324; shift_adder #(17, 11, 1, 1, 18, 6, 0) op_2324 (v335[16:0], v672[10:0], v2324[17:0]); // 2.0
    wire [17:0] v2325; shift_adder #(11, 17, 1, 1, 18, -6, 0) op_2325 (v367[10:0], v677[16:0], v2325[17:0]); // 2.0
    wire [21:0] v2326; shift_adder #(12, 21, 1, 1, 22, -10, 0) op_2326 (v383[11:0], v624[20:0], v2326[21:0]); // 2.0
    wire [13:0] v2327; shift_adder #(12, 10, 1, 1, 14, 4, 0) op_2327 (v174[11:0], v254[9:0], v2327[13:0]); // 2.0
    wire [16:0] v2328; shift_adder #(11, 17, 1, 1, 17, -4, 0) op_2328 (v577[10:0], v306[16:0], v2328[16:0]); // 2.0
    wire [32:0] v2329; shift_adder #(14, 33, 1, 1, 33, -16, 0) op_2329 (v571[13:0], v726[32:0], v2329[32:0]); // 2.0
    wire [11:0] v2330; shift_adder #(11, 11, 1, 1, 12, 0, 0) op_2330 (v162[10:0], v154[10:0], v2330[11:0]); // 2.0
    wire [13:0] v2331; shift_adder #(12, 14, 1, 1, 14, 0, 0) op_2331 (v227[11:0], v454[13:0], v2331[13:0]); // 2.0
    wire [37:0] v2332; shift_adder #(12, 8, 1, 1, 38, 29, 1) op_2332 (v579[11:0], v93[7:0], v2332[37:0]); // 2.0
    wire [12:0] v2333; shift_adder #(13, 10, 1, 1, 13, 0, 0) op_2333 (v601[12:0], v727[9:0], v2333[12:0]); // 2.0
    wire [11:0] v2334; shift_adder #(8, 11, 1, 1, 12, -2, 0) op_2334 (v93[7:0], v393[10:0], v2334[11:0]); // 2.0
    wire [10:0] v2335; shift_adder #(11, 9, 1, 1, 11, 0, 0) op_2335 (v728[10:0], v302[8:0], v2335[10:0]); // 2.0
    wire [14:0] v2336; shift_adder #(14, 12, 1, 1, 15, -1, 0) op_2336 (v499[13:0], v383[11:0], v2336[14:0]); // 2.0
    wire [11:0] v2337; shift_adder #(12, 10, 1, 1, 12, 1, 0) op_2337 (v457[11:0], v722[9:0], v2337[11:0]); // 2.0
    wire [11:0] v2338; shift_adder #(11, 11, 1, 1, 12, 1, 0) op_2338 (v622[10:0], v729[10:0], v2338[11:0]); // 2.0
    wire [9:0] v2339; shift_adder #(8, 9, 1, 1, 10, 0, 0) op_2339 (v126[7:0], v477[8:0], v2339[9:0]); // 2.0
    wire [11:0] v2340; shift_adder #(11, 11, 1, 1, 12, -1, 0) op_2340 (v206[10:0], v294[10:0], v2340[11:0]); // 2.0
    wire [11:0] v2341; shift_adder #(8, 11, 1, 1, 12, -3, 1) op_2341 (v68[7:0], v319[10:0], v2341[11:0]); // 2.0
    wire [38:0] v2342; shift_adder #(10, 15, 1, 1, 39, -29, 1) op_2342 (v489[9:0], v308[14:0], v2342[38:0]); // 2.0
    wire [29:0] v2343; shift_adder #(12, 14, 1, 1, 30, 16, 1) op_2343 (v174[11:0], v481[13:0], v2343[29:0]); // 2.0
    wire [25:0] v2344; shift_adder #(25, 11, 1, 1, 26, 15, 0) op_2344 (v537[24:0], v338[10:0], v2344[25:0]); // 2.0
    wire [16:0] v2345; shift_adder #(9, 10, 1, 1, 17, -7, 0) op_2345 (v369[8:0], v252[9:0], v2345[16:0]); // 2.0
    wire [10:0] v2346; shift_adder #(8, 11, 1, 1, 11, 0, 0) op_2346 (v82[7:0], v294[10:0], v2346[10:0]); // 2.0
    wire [25:0] v2347; shift_adder #(11, 11, 1, 1, 26, 15, 0) op_2347 (v362[10:0], v242[10:0], v2347[25:0]); // 2.0
    wire [11:0] v2348; shift_adder #(12, 10, 1, 1, 12, 1, 0) op_2348 (v137[11:0], v254[9:0], v2348[11:0]); // 2.0
    wire [21:0] v2349; shift_adder #(8, 11, 1, 1, 22, -13, 0) op_2349 (v102[7:0], v201[10:0], v2349[21:0]); // 2.0
    wire [12:0] v2350; shift_adder #(13, 11, 1, 1, 13, 1, 0) op_2350 (v449[12:0], v163[10:0], v2350[12:0]); // 2.0
    wire [19:0] v2351; shift_adder #(13, 10, 1, 1, 20, 10, 0) op_2351 (v573[12:0], v569[9:0], v2351[19:0]); // 2.0
    wire [11:0] v2352; shift_adder #(11, 11, 1, 1, 12, 1, 0) op_2352 (v169[10:0], v218[10:0], v2352[11:0]); // 2.0
    wire [12:0] v2353; shift_adder #(12, 12, 1, 1, 13, 0, 1) op_2353 (v285[11:0], v388[11:0], v2353[12:0]); // 2.0
    wire [12:0] v2354; shift_adder #(11, 10, 1, 1, 13, 2, 0) op_2354 (v361[10:0], v282[9:0], v2354[12:0]); // 2.0
    wire [21:0] v2355; shift_adder #(11, 21, 1, 1, 22, -10, 0) op_2355 (v141[10:0], v624[20:0], v2355[21:0]); // 2.0
    wire [13:0] v2356; shift_adder #(10, 13, 1, 1, 14, -3, 0) op_2356 (v263[9:0], v346[12:0], v2356[13:0]); // 2.0
    wire [14:0] v2357; shift_adder #(15, 11, 1, 1, 15, 1, 0) op_2357 (v313[14:0], v237[10:0], v2357[14:0]); // 2.0
    wire [12:0] v2358; shift_adder #(12, 11, 1, 1, 13, -1, 0) op_2358 (v227[11:0], v155[10:0], v2358[12:0]); // 2.0
    wire [26:0] v2359; shift_adder #(11, 11, 1, 1, 27, -16, 0) op_2359 (v294[10:0], v317[10:0], v2359[26:0]); // 2.0
    wire [17:0] v2360; shift_adder #(10, 16, 1, 1, 18, -7, 0) op_2360 (v730[9:0], v731[15:0], v2360[17:0]); // 2.0
    wire [24:0] v2361; shift_adder #(8, 10, 1, 1, 25, -16, 1) op_2361 (v87[7:0], v282[9:0], v2361[24:0]); // 2.0
    wire [15:0] v2362; shift_adder #(11, 13, 1, 1, 16, -5, 0) op_2362 (v602[10:0], v506[12:0], v2362[15:0]); // 2.0
    wire [13:0] v2363; shift_adder #(11, 11, 1, 1, 14, 3, 0) op_2363 (v277[10:0], v518[10:0], v2363[13:0]); // 2.0
    wire [13:0] v2364; shift_adder #(11, 9, 1, 1, 14, 4, 0) op_2364 (v212[10:0], v384[8:0], v2364[13:0]); // 2.0
    wire [32:0] v2365; shift_adder #(11, 13, 1, 1, 33, -22, 1) op_2365 (v157[10:0], v449[12:0], v2365[32:0]); // 2.0
    wire [18:0] v2366; shift_adder #(11, 19, 1, 1, 19, -4, 0) op_2366 (v177[10:0], v732[18:0], v2366[18:0]); // 2.0
    wire [11:0] v2367; shift_adder #(12, 11, 1, 1, 12, 0, 0) op_2367 (v404[11:0], v418[10:0], v2367[11:0]); // 2.0
    wire [14:0] v2368; shift_adder #(11, 11, 1, 1, 15, 4, 0) op_2368 (v134[10:0], v714[10:0], v2368[14:0]); // 2.0
    wire [12:0] v2369; shift_adder #(9, 12, 1, 1, 13, -2, 0) op_2369 (v403[8:0], v734[11:0], v2369[12:0]); // 2.0
    wire [12:0] v2370; shift_adder #(12, 12, 1, 1, 13, 0, 0) op_2370 (v550[11:0], v553[11:0], v2370[12:0]); // 2.0
    wire [12:0] v2371; shift_adder #(8, 11, 1, 1, 13, -4, 1) op_2371 (v84[7:0], v177[10:0], v2371[12:0]); // 2.0
    wire [11:0] v2372; shift_adder #(11, 11, 1, 1, 12, 0, 0) op_2372 (v497[10:0], v141[10:0], v2372[11:0]); // 2.0
    wire [16:0] v2373; shift_adder #(17, 13, 1, 1, 17, 3, 0) op_2373 (v689[16:0], v735[12:0], v2373[16:0]); // 2.0
    wire [11:0] v2374; shift_adder #(12, 11, 1, 1, 12, 0, 0) op_2374 (v180[11:0], v277[10:0], v2374[11:0]); // 2.0
    wire [12:0] v2375; shift_adder #(11, 11, 1, 1, 13, 2, 1) op_2375 (v140[10:0], v234[10:0], v2375[12:0]); // 2.0
    wire [12:0] v2376; shift_adder #(12, 11, 1, 1, 13, -1, 0) op_2376 (v267[11:0], v424[10:0], v2376[12:0]); // 2.0
    wire [11:0] v2377; shift_adder #(11, 11, 1, 1, 12, -1, 0) op_2377 (v420[10:0], v172[10:0], v2377[11:0]); // 2.0
    wire [11:0] v2378; shift_adder #(11, 9, 1, 1, 12, -1, 0) op_2378 (v736[10:0], v220[8:0], v2378[11:0]); // 2.0
    wire [13:0] v2379; shift_adder #(11, 12, 1, 1, 14, 2, 0) op_2379 (v197[10:0], v146[11:0], v2379[13:0]); // 2.0
    wire [16:0] v2380; shift_adder #(14, 15, 1, 1, 17, -3, 0) op_2380 (v444[13:0], v253[14:0], v2380[16:0]); // 2.0
    wire [14:0] v2381; shift_adder #(11, 11, 1, 1, 15, 4, 0) op_2381 (v418[10:0], v211[10:0], v2381[14:0]); // 2.0
    wire [11:0] v2382; shift_adder #(11, 11, 1, 1, 12, 0, 0) op_2382 (v300[10:0], v329[10:0], v2382[11:0]); // 2.0
    wire [14:0] v2383; shift_adder #(12, 15, 1, 1, 15, -2, 0) op_2383 (v280[11:0], v649[14:0], v2383[14:0]); // 2.0
    wire [19:0] v2384; shift_adder #(20, 12, 1, 1, 20, 7, 0) op_2384 (v737[19:0], v265[11:0], v2384[19:0]); // 2.0
    wire [11:0] v2385; shift_adder #(11, 11, 1, 1, 12, 0, 0) op_2385 (v738[10:0], v367[10:0], v2385[11:0]); // 2.0
    wire [12:0] v2386; shift_adder #(12, 12, 1, 1, 13, 1, 0) op_2386 (v447[11:0], v398[11:0], v2386[12:0]); // 2.0
    wire [13:0] v2387; shift_adder #(12, 11, 1, 1, 14, 3, 0) op_2387 (v325[11:0], v238[10:0], v2387[13:0]); // 2.0
    wire [11:0] v2388; shift_adder #(10, 11, 1, 1, 12, -1, 0) op_2388 (v739[9:0], v659[10:0], v2388[11:0]); // 2.0
    wire [17:0] v2389; shift_adder #(16, 9, 1, 1, 18, 8, 0) op_2389 (v426[15:0], v441[8:0], v2389[17:0]); // 2.0
    wire [12:0] v2390; shift_adder #(11, 10, 1, 1, 13, 3, 1) op_2390 (v177[10:0], v248[9:0], v2390[12:0]); // 2.0
    wire [14:0] v2391; shift_adder #(14, 10, 1, 1, 15, 4, 0) op_2391 (v603[13:0], v130[9:0], v2391[14:0]); // 2.0
    wire [12:0] v2392; shift_adder #(11, 12, 1, 1, 13, -1, 0) op_2392 (v136[10:0], v462[11:0], v2392[12:0]); // 2.0
    wire [11:0] v2393; shift_adder #(10, 11, 1, 1, 12, -1, 0) op_2393 (v225[9:0], v287[10:0], v2393[11:0]); // 2.0
    wire [35:0] v2394; shift_adder #(11, 8, 1, 1, 36, 27, 1) op_2394 (v208[10:0], v109[7:0], v2394[35:0]); // 2.0
    wire [12:0] v2395; shift_adder #(11, 11, 1, 1, 13, 2, 0) op_2395 (v201[10:0], v430[10:0], v2395[12:0]); // 2.0
    wire [13:0] v2396; shift_adder #(10, 11, 1, 1, 14, -4, 0) op_2396 (v466[9:0], v740[10:0], v2396[13:0]); // 2.0
    wire [16:0] v2397; shift_adder #(11, 12, 1, 1, 17, 5, 1) op_2397 (v158[10:0], v404[11:0], v2397[16:0]); // 2.0
    wire [19:0] v2398; shift_adder #(10, 18, 1, 1, 20, -10, 0) op_2398 (v366[9:0], v741[17:0], v2398[19:0]); // 2.0
    wire [11:0] v2399; shift_adder #(11, 11, 1, 1, 12, -1, 0) op_2399 (v139[10:0], v312[10:0], v2399[11:0]); // 2.0
    wire [12:0] v2400; shift_adder #(12, 11, 1, 1, 13, 1, 0) op_2400 (v389[11:0], v396[10:0], v2400[12:0]); // 2.0
    wire [10:0] v2401; shift_adder #(11, 9, 1, 1, 11, 0, 0) op_2401 (v659[10:0], v351[8:0], v2401[10:0]); // 2.0
    wire [11:0] v2402; shift_adder #(11, 11, 1, 1, 12, 0, 0) op_2402 (v328[10:0], v218[10:0], v2402[11:0]); // 2.0
    wire [22:0] v2403; shift_adder #(23, 12, 1, 1, 23, 9, 0) op_2403 (v440[22:0], v280[11:0], v2403[22:0]); // 2.0
    wire [11:0] v2404; shift_adder #(11, 9, 1, 1, 12, 1, 0) op_2404 (v241[10:0], v490[8:0], v2404[11:0]); // 2.0
    wire [11:0] v2405; shift_adder #(11, 11, 1, 1, 12, -1, 0) op_2405 (v144[10:0], v284[10:0], v2405[11:0]); // 2.0
    wire [16:0] v2406; shift_adder #(16, 16, 1, 1, 17, 0, 0) op_2406 (v731[15:0], v240[15:0], v2406[16:0]); // 2.0
    wire [12:0] v2407; shift_adder #(13, 10, 1, 1, 13, 2, 0) op_2407 (v742[12:0], v678[9:0], v2407[12:0]); // 2.0
    wire [24:0] v2408; shift_adder #(11, 25, 1, 1, 25, -11, 0) op_2408 (v201[10:0], v595[24:0], v2408[24:0]); // 2.0
    wire [13:0] v2409; shift_adder #(13, 9, 1, 1, 14, 4, 0) op_2409 (v598[12:0], v138[8:0], v2409[13:0]); // 2.0
    wire [11:0] v2410; shift_adder #(11, 11, 1, 1, 12, 1, 0) op_2410 (v234[10:0], v270[10:0], v2410[11:0]); // 2.0
    wire [10:0] v2411; shift_adder #(10, 11, 1, 1, 11, 0, 0) op_2411 (v282[9:0], v176[10:0], v2411[10:0]); // 2.0
    wire [13:0] v2412; shift_adder #(11, 11, 1, 1, 14, -3, 1) op_2412 (v255[10:0], v352[10:0], v2412[13:0]); // 2.0
    wire [15:0] v2413; shift_adder #(11, 15, 1, 1, 16, -4, 0) op_2413 (v361[10:0], v630[14:0], v2413[15:0]); // 2.0
    wire [14:0] v2414; shift_adder #(11, 11, 1, 1, 15, -4, 1) op_2414 (v219[10:0], v208[10:0], v2414[14:0]); // 2.0
    wire [21:0] v2415; shift_adder #(18, 22, 1, 1, 22, 0, 0) op_2415 (v535[17:0], v743[21:0], v2415[21:0]); // 2.0
    wire [11:0] v2416; shift_adder #(12, 11, 1, 1, 12, 0, 0) op_2416 (v325[11:0], v245[10:0], v2416[11:0]); // 2.0
    wire [13:0] v2417; shift_adder #(13, 13, 1, 1, 14, 0, 0) op_2417 (v601[12:0], v744[12:0], v2417[13:0]); // 2.0
    wire [11:0] v2418; shift_adder #(11, 11, 1, 1, 12, 0, 0) op_2418 (v185[10:0], v714[10:0], v2418[11:0]); // 2.0
    wire [13:0] v2419; shift_adder #(11, 11, 1, 1, 14, 3, 0) op_2419 (v745[10:0], v478[10:0], v2419[13:0]); // 2.0
    wire [15:0] v2420; shift_adder #(13, 10, 1, 1, 16, 6, 0) op_2420 (v344[12:0], v746[9:0], v2420[15:0]); // 2.0
    wire [12:0] v2421; shift_adder #(11, 11, 1, 1, 13, 2, 0) op_2421 (v145[10:0], v217[10:0], v2421[12:0]); // 2.0
    wire [11:0] v2422; shift_adder #(11, 11, 1, 1, 12, -1, 0) op_2422 (v747[10:0], v179[10:0], v2422[11:0]); // 2.0
    wire [12:0] v2423; shift_adder #(12, 9, 1, 1, 13, 3, 0) op_2423 (v389[11:0], v479[8:0], v2423[12:0]); // 2.0
    wire [11:0] v2424; shift_adder #(11, 11, 1, 1, 12, -1, 0) op_2424 (v148[10:0], v298[10:0], v2424[11:0]); // 2.0
    wire [11:0] v2425; shift_adder #(11, 11, 1, 1, 12, -1, 0) op_2425 (v175[10:0], v319[10:0], v2425[11:0]); // 2.0
    wire [10:0] v2426; shift_adder #(9, 11, 1, 1, 11, 0, 0) op_2426 (v490[8:0], v250[10:0], v2426[10:0]); // 2.0
    wire [39:0] v2427; shift_adder #(10, 12, 1, 1, 40, -30, 1) op_2427 (v748[9:0], v523[11:0], v2427[39:0]); // 2.0
    wire [10:0] v2428; shift_adder #(11, 9, 1, 1, 11, 0, 0) op_2428 (v329[10:0], v556[8:0], v2428[10:0]); // 2.0
    wire [11:0] v2429; shift_adder #(10, 11, 1, 1, 12, -1, 0) op_2429 (v585[9:0], v386[10:0], v2429[11:0]); // 2.0
    wire [13:0] v2430; shift_adder #(11, 13, 1, 1, 14, -3, 0) op_2430 (v393[10:0], v573[12:0], v2430[13:0]); // 2.0
    wire [10:0] v2431; shift_adder #(9, 10, 1, 1, 11, 0, 0) op_2431 (v302[8:0], v705[9:0], v2431[10:0]); // 2.0
    wire [14:0] v2432; shift_adder #(12, 14, 1, 1, 15, -2, 0) op_2432 (v523[11:0], v603[13:0], v2432[14:0]); // 2.0
    wire [13:0] v2433; shift_adder #(9, 14, 1, 1, 14, -3, 0) op_2433 (v749[8:0], v412[13:0], v2433[13:0]); // 2.0
    wire [11:0] v2434; shift_adder #(10, 11, 1, 1, 12, -1, 0) op_2434 (v469[9:0], v379[10:0], v2434[11:0]); // 2.0
    wire [23:0] v2435; shift_adder #(11, 24, 1, 1, 24, -11, 0) op_2435 (v328[10:0], v559[23:0], v2435[23:0]); // 2.0
    wire [12:0] v2436; shift_adder #(11, 10, 1, 1, 13, 3, 0) op_2436 (v750[10:0], v254[9:0], v2436[12:0]); // 2.0
    wire [12:0] v2437; shift_adder #(12, 12, 1, 1, 13, 1, 0) op_2437 (v202[11:0], v347[11:0], v2437[12:0]); // 2.0
    wire [13:0] v2438; shift_adder #(12, 12, 1, 1, 14, -2, 0) op_2438 (v464[11:0], v207[11:0], v2438[13:0]); // 2.0
    wire [17:0] v2439; shift_adder #(17, 10, 1, 1, 18, 8, 0) op_2439 (v751[16:0], v632[9:0], v2439[17:0]); // 2.0
    wire [14:0] v2440; shift_adder #(11, 12, 1, 1, 15, 3, 0) op_2440 (v246[10:0], v532[11:0], v2440[14:0]); // 2.0
    wire [12:0] v2441; shift_adder #(12, 12, 1, 1, 13, 1, 0) op_2441 (v586[11:0], v174[11:0], v2441[12:0]); // 2.0
    wire [12:0] v2442; shift_adder #(11, 12, 1, 1, 13, -2, 0) op_2442 (v752[10:0], v279[11:0], v2442[12:0]); // 2.0
    wire [9:0] v2443; shift_adder #(9, 9, 1, 1, 10, 0, 0) op_2443 (v479[8:0], v128[8:0], v2443[9:0]); // 2.0
    wire [12:0] v2444; shift_adder #(11, 12, 1, 1, 13, 1, 0) op_2444 (v266[10:0], v532[11:0], v2444[12:0]); // 2.0
    wire [19:0] v2445; shift_adder #(9, 19, 1, 1, 20, -10, 0) op_2445 (v490[8:0], v376[18:0], v2445[19:0]); // 2.0
    wire [12:0] v2446; shift_adder #(11, 10, 1, 1, 13, 3, 0) op_2446 (v362[10:0], v421[9:0], v2446[12:0]); // 2.0
    wire [11:0] v2447; shift_adder #(9, 11, 1, 1, 12, -2, 0) op_2447 (v369[8:0], v219[10:0], v2447[11:0]); // 2.0
    wire [18:0] v2448; shift_adder #(11, 19, 1, 1, 19, -6, 0) op_2448 (v487[10:0], v558[18:0], v2448[18:0]); // 2.0
    wire [15:0] v2449; shift_adder #(15, 11, 1, 1, 16, 4, 0) op_2449 (v295[14:0], v162[10:0], v2449[15:0]); // 2.0
    wire [12:0] v2450; shift_adder #(11, 12, 1, 1, 13, 1, 0) op_2450 (v276[10:0], v137[11:0], v2450[12:0]); // 2.0
    wire [22:0] v2451; shift_adder #(12, 23, 1, 1, 23, -10, 0) op_2451 (v657[11:0], v753[22:0], v2451[22:0]); // 2.0
    wire [13:0] v2452; shift_adder #(11, 13, 1, 1, 14, -2, 0) op_2452 (v396[10:0], v344[12:0], v2452[13:0]); // 2.0
    wire [18:0] v2453; shift_adder #(18, 17, 1, 1, 19, 2, 0) op_2453 (v493[17:0], v689[16:0], v2453[18:0]); // 2.0
    wire [35:0] v2454; shift_adder #(11, 11, 1, 1, 36, -25, 1) op_2454 (v134[10:0], v269[10:0], v2454[35:0]); // 2.0
    wire [11:0] v2455; shift_adder #(11, 11, 1, 1, 12, -1, 0) op_2455 (v377[10:0], v155[10:0], v2455[11:0]); // 2.0
    wire [12:0] v2456; shift_adder #(9, 11, 1, 1, 13, -3, 0) op_2456 (v395[8:0], v135[10:0], v2456[12:0]); // 2.0
    wire [13:0] v2457; shift_adder #(13, 9, 1, 1, 14, 3, 0) op_2457 (v189[12:0], v754[8:0], v2457[13:0]); // 2.0
    wire [16:0] v2458; shift_adder #(15, 13, 1, 1, 17, -2, 0) op_2458 (v482[14:0], v755[12:0], v2458[16:0]); // 2.0
    wire [10:0] v2459; shift_adder #(11, 10, 1, 1, 11, 0, 0) op_2459 (v430[10:0], v549[9:0], v2459[10:0]); // 2.0
    wire [21:0] v2460; shift_adder #(11, 11, 1, 1, 22, 11, 1) op_2460 (v163[10:0], v361[10:0], v2460[21:0]); // 2.0
    wire [13:0] v2461; shift_adder #(12, 11, 1, 1, 14, -2, 0) op_2461 (v495[11:0], v145[10:0], v2461[13:0]); // 2.0
    wire [12:0] v2462; shift_adder #(12, 12, 1, 1, 13, -1, 0) op_2462 (v453[11:0], v257[11:0], v2462[12:0]); // 2.0
    wire [16:0] v2463; shift_adder #(8, 11, 1, 1, 17, 6, 0) op_2463 (v96[7:0], v168[10:0], v2463[16:0]); // 2.0
    wire [12:0] v2464; shift_adder #(10, 11, 1, 1, 13, -3, 0) op_2464 (v463[9:0], v756[10:0], v2464[12:0]); // 2.0
    wire [17:0] v2465; shift_adder #(12, 17, 1, 1, 18, 1, 0) op_2465 (v589[11:0], v757[16:0], v2465[17:0]); // 2.0
    wire [14:0] v2466; shift_adder #(12, 10, 1, 1, 15, 5, 0) op_2466 (v407[11:0], v510[9:0], v2466[14:0]); // 2.0
    wire [10:0] v2467; shift_adder #(9, 9, 1, 1, 11, 1, 0) op_2467 (v758[8:0], v128[8:0], v2467[10:0]); // 2.0
    wire [16:0] v2468; shift_adder #(17, 11, 1, 1, 17, 4, 0) op_2468 (v759[16:0], v343[10:0], v2468[16:0]); // 2.0
    wire [12:0] v2469; shift_adder #(11, 11, 1, 1, 13, 2, 0) op_2469 (v298[10:0], v216[10:0], v2469[12:0]); // 2.0
    wire [18:0] v2470; shift_adder #(13, 18, 1, 1, 19, -5, 0) op_2470 (v296[12:0], v167[17:0], v2470[18:0]); // 2.0
    wire [11:0] v2471; shift_adder #(11, 11, 1, 1, 12, 1, 0) op_2471 (v223[10:0], v329[10:0], v2471[11:0]); // 2.0
    wire [10:0] v2472; shift_adder #(9, 11, 1, 1, 11, 0, 0) op_2472 (v220[8:0], v212[10:0], v2472[10:0]); // 2.0
    wire [11:0] v2473; shift_adder #(11, 11, 1, 1, 12, 0, 0) op_2473 (v367[10:0], v178[10:0], v2473[11:0]); // 2.0
    wire [17:0] v2474; shift_adder #(12, 12, 1, 1, 18, -6, 1) op_2474 (v398[11:0], v398[11:0], v2474[17:0]); // 2.0
    wire [20:0] v2475; shift_adder #(11, 21, 1, 1, 21, -6, 0) op_2475 (v190[10:0], v760[20:0], v2475[20:0]); // 2.0
    wire [37:0] v2476; shift_adder #(9, 38, 1, 1, 38, -28, 0) op_2476 (v360[8:0], v761[37:0], v2476[37:0]); // 2.0
    wire [33:0] v2477; shift_adder #(11, 11, 1, 1, 34, -23, 1) op_2477 (v268[10:0], v379[10:0], v2477[33:0]); // 2.0
    wire [11:0] v2478; shift_adder #(10, 9, 1, 1, 12, 2, 0) op_2478 (v307[9:0], v538[8:0], v2478[11:0]); // 2.0
    wire [16:0] v2479; shift_adder #(17, 14, 1, 1, 17, 1, 0) op_2479 (v533[16:0], v555[13:0], v2479[16:0]); // 2.0
    wire [28:0] v2480; shift_adder #(9, 29, 1, 1, 29, -19, 0) op_2480 (v405[8:0], v439[28:0], v2480[28:0]); // 2.0
    wire [11:0] v2481; shift_adder #(12, 11, 1, 1, 12, 0, 0) op_2481 (v500[11:0], v275[10:0], v2481[11:0]); // 2.0
    wire [13:0] v2482; shift_adder #(11, 12, 1, 1, 14, -3, 0) op_2482 (v217[10:0], v762[11:0], v2482[13:0]); // 2.0
    wire [15:0] v2483; shift_adder #(11, 15, 1, 1, 16, -5, 0) op_2483 (v168[10:0], v313[14:0], v2483[15:0]); // 2.0
    wire [18:0] v2484; shift_adder #(19, 10, 1, 1, 19, 6, 0) op_2484 (v539[18:0], v763[9:0], v2484[18:0]); // 2.0
    wire [19:0] v2485; shift_adder #(20, 12, 1, 1, 20, 7, 0) op_2485 (v764[19:0], v137[11:0], v2485[19:0]); // 2.0
    wire [12:0] v2486; shift_adder #(9, 12, 1, 1, 13, -3, 0) op_2486 (v351[8:0], v397[11:0], v2486[12:0]); // 2.0
    wire [12:0] v2487; shift_adder #(12, 11, 1, 1, 13, 1, 0) op_2487 (v657[11:0], v213[10:0], v2487[12:0]); // 2.0
    wire [19:0] v2488; shift_adder #(19, 14, 1, 1, 20, 6, 0) op_2488 (v536[18:0], v765[13:0], v2488[19:0]); // 2.0
    wire [26:0] v2489; shift_adder #(23, 12, 1, 1, 27, 15, 0) op_2489 (v766[22:0], v204[11:0], v2489[26:0]); // 2.0
    wire [18:0] v2490; shift_adder #(12, 18, 1, 1, 19, -7, 0) op_2490 (v507[11:0], v633[17:0], v2490[18:0]); // 2.0
    wire [11:0] v2491; shift_adder #(12, 11, 1, 1, 12, 0, 0) op_2491 (v183[11:0], v277[10:0], v2491[11:0]); // 2.0
    wire [14:0] v2492; shift_adder #(14, 13, 1, 1, 15, 1, 0) op_2492 (v460[13:0], v451[12:0], v2492[14:0]); // 2.0
    wire [18:0] v2493; shift_adder #(19, 11, 1, 1, 19, 6, 0) op_2493 (v376[18:0], v147[10:0], v2493[18:0]); // 2.0
    wire [12:0] v2494; shift_adder #(13, 11, 1, 1, 13, 1, 0) op_2494 (v359[12:0], v277[10:0], v2494[12:0]); // 2.0
    wire [11:0] v2495; shift_adder #(11, 11, 1, 1, 12, -1, 0) op_2495 (v289[10:0], v156[10:0], v2495[11:0]); // 2.0
    wire [13:0] v2496; shift_adder #(12, 13, 1, 1, 14, 1, 0) op_2496 (v397[11:0], v578[12:0], v2496[13:0]); // 2.0
    wire [16:0] v2497; shift_adder #(14, 16, 1, 1, 17, -3, 0) op_2497 (v499[13:0], v426[15:0], v2497[16:0]); // 2.0
    wire [14:0] v2498; shift_adder #(13, 10, 1, 1, 15, 4, 0) op_2498 (v346[12:0], v584[9:0], v2498[14:0]); // 2.0
    wire [12:0] v2499; shift_adder #(11, 13, 1, 1, 13, 0, 0) op_2499 (v206[10:0], v625[12:0], v2499[12:0]); // 2.0
    wire [14:0] v2500; shift_adder #(12, 15, 1, 1, 15, -1, 0) op_2500 (v292[11:0], v767[14:0], v2500[14:0]); // 2.0
    wire [12:0] v2501; shift_adder #(12, 11, 1, 1, 13, 1, 0) op_2501 (v550[11:0], v185[10:0], v2501[12:0]); // 2.0
    wire [11:0] v2502; shift_adder #(11, 11, 1, 1, 12, 0, 0) op_2502 (v400[10:0], v175[10:0], v2502[11:0]); // 2.0
    wire [13:0] v2503; shift_adder #(13, 11, 1, 1, 14, 2, 0) op_2503 (v601[12:0], v145[10:0], v2503[13:0]); // 2.0
    wire [34:0] v2504; shift_adder #(12, 11, 1, 1, 35, -23, 1) op_2504 (v355[11:0], v768[10:0], v2504[34:0]); // 2.0
    wire [16:0] v2505; shift_adder #(14, 16, 1, 1, 17, -3, 0) op_2505 (v590[13:0], v426[15:0], v2505[16:0]); // 2.0
    wire [11:0] v2506; shift_adder #(11, 11, 1, 1, 12, 1, 0) op_2506 (v181[10:0], v769[10:0], v2506[11:0]); // 2.0
    wire [22:0] v2507; shift_adder #(11, 22, 1, 1, 23, -12, 0) op_2507 (v269[10:0], v371[21:0], v2507[22:0]); // 2.0
    wire [28:0] v2508; shift_adder #(11, 28, 1, 1, 29, -17, 0) op_2508 (v145[10:0], v593[27:0], v2508[28:0]); // 2.0
    wire [13:0] v2509; shift_adder #(14, 11, 1, 1, 14, 2, 0) op_2509 (v226[13:0], v300[10:0], v2509[13:0]); // 2.0
    wire [13:0] v2510; shift_adder #(12, 10, 1, 1, 14, 4, 0) op_2510 (v337[11:0], v273[9:0], v2510[13:0]); // 2.0
    wire [13:0] v2511; shift_adder #(11, 11, 1, 1, 14, -3, 0) op_2511 (v379[10:0], v132[10:0], v2511[13:0]); // 2.0
    wire [18:0] v2512; shift_adder #(18, 13, 1, 1, 19, 6, 0) op_2512 (v770[17:0], v771[12:0], v2512[18:0]); // 3.0
    wire [15:0] v2513; shift_adder #(11, 11, 1, 1, 16, -5, 0) op_2513 (v131[10:0], v772[10:0], v2513[15:0]); // 3.0
    wire [23:0] v2514; shift_adder #(11, 17, 1, 1, 24, -13, 0) op_2514 (v133[10:0], v773[16:0], v2514[23:0]); // 3.0
    wire [21:0] v2515; shift_adder #(22, 12, 1, 1, 22, 9, 0) op_2515 (v774[21:0], v775[11:0], v2515[21:0]); // 3.0
    wire [18:0] v2516; shift_adder #(11, 19, 1, 1, 19, -2, 0) op_2516 (v140[10:0], v776[18:0], v2516[18:0]); // 3.0
    wire [21:0] v2517; shift_adder #(21, 16, 1, 1, 22, 6, 0) op_2517 (v777[20:0], v778[15:0], v2517[21:0]); // 3.0
    wire [21:0] v2518; shift_adder #(12, 15, 1, 1, 22, -10, 1) op_2518 (v146[11:0], v779[14:0], v2518[21:0]); // 3.0
    wire [23:0] v2519; shift_adder #(13, 24, 1, 1, 24, -2, 1) op_2519 (v149[12:0], v780[23:0], v2519[23:0]); // 3.0
    wire [25:0] v2520; shift_adder #(12, 19, 1, 1, 26, 7, 0) op_2520 (v137[11:0], v782[18:0], v2520[25:0]); // 3.0
    wire [24:0] v2521; shift_adder #(17, 25, 1, 1, 25, -7, 0) op_2521 (v783[16:0], v784[24:0], v2521[24:0]); // 3.0
    wire [12:0] v2522; shift_adder #(11, 11, 1, 1, 13, 1, 1) op_2522 (v161[10:0], v785[10:0], v2522[12:0]); // 3.0
    wire [14:0] v2523; shift_adder #(14, 14, 1, 1, 15, 0, 0) op_2523 (v786[13:0], v787[13:0], v2523[14:0]); // 3.0
    wire [24:0] v2524; shift_adder #(23, 18, 1, 1, 25, 7, 0) op_2524 (v788[22:0], v789[17:0], v2524[24:0]); // 3.0
    wire [27:0] v2525; shift_adder #(11, 25, 1, 1, 28, 3, 1) op_2525 (v145[10:0], v791[24:0], v2525[27:0]); // 3.0
    wire [13:0] v2526; shift_adder #(8, 13, 1, 1, 14, 1, 0) op_2526 (v92[7:0], v792[12:0], v2526[13:0]); // 3.0
    wire [23:0] v2527; shift_adder #(12, 13, 1, 1, 24, -12, 0) op_2527 (v174[11:0], v793[12:0], v2527[23:0]); // 3.0
    wire [12:0] v2528; shift_adder #(11, 12, 1, 1, 13, -1, 0) op_2528 (v176[10:0], v794[11:0], v2528[12:0]); // 3.0
    wire [16:0] v2529; shift_adder #(8, 13, 1, 1, 17, -8, 1) op_2529 (v112[7:0], v795[12:0], v2529[16:0]); // 3.0
    wire [22:0] v2530; shift_adder #(8, 12, 1, 1, 23, 11, 1) op_2530 (v92[7:0], v797[11:0], v2530[22:0]); // 3.0
    wire [27:0] v2531; shift_adder #(27, 14, 1, 1, 28, 14, 0) op_2531 (v798[26:0], v799[13:0], v2531[27:0]); // 3.0
    wire [13:0] v2532; shift_adder #(13, 12, 1, 1, 14, -1, 0) op_2532 (v800[12:0], v801[11:0], v2532[13:0]); // 3.0
    wire [26:0] v2533; shift_adder #(13, 26, 1, 1, 27, -13, 0) op_2533 (v189[12:0], v802[25:0], v2533[26:0]); // 3.0
    wire [13:0] v2534; shift_adder #(13, 13, 1, 1, 14, 0, 1) op_2534 (v192[12:0], v803[12:0], v2534[13:0]); // 3.0
    wire [21:0] v2535; shift_adder #(22, 19, 1, 1, 22, 0, 0) op_2535 (v804[21:0], v805[18:0], v2535[21:0]); // 3.0
    wire [20:0] v2536; shift_adder #(20, 14, 1, 1, 21, 7, 0) op_2536 (v806[19:0], v807[13:0], v2536[20:0]); // 3.0
    wire [12:0] v2537; shift_adder #(11, 12, 1, 1, 13, 0, 1) op_2537 (v199[10:0], v808[11:0], v2537[12:0]); // 3.0
    wire [26:0] v2538; shift_adder #(8, 20, 1, 1, 27, 7, 0) op_2538 (v118[7:0], v809[19:0], v2538[26:0]); // 3.0
    wire [30:0] v2539; shift_adder #(8, 26, 1, 1, 31, -22, 0) op_2539 (v110[7:0], v810[25:0], v2539[30:0]); // 3.0
    wire [30:0] v2540; shift_adder #(23, 29, 1, 1, 31, -8, 0) op_2540 (v811[22:0], v812[28:0], v2540[30:0]); // 3.0
    wire [16:0] v2541; shift_adder #(13, 16, 1, 1, 17, -3, 0) op_2541 (v813[12:0], v814[15:0], v2541[16:0]); // 3.0
    wire [17:0] v2542; shift_adder #(15, 18, 1, 1, 18, -1, 0) op_2542 (v815[14:0], v816[17:0], v2542[17:0]); // 3.0
    wire [17:0] v2543; shift_adder #(13, 13, 1, 1, 18, -5, 0) op_2543 (v817[12:0], v818[12:0], v2543[17:0]); // 3.0
    wire [18:0] v2544; shift_adder #(11, 17, 1, 1, 19, -8, 0) op_2544 (v215[10:0], v819[16:0], v2544[18:0]); // 3.0
    wire [12:0] v2545; shift_adder #(12, 9, 1, 1, 13, 2, 0) op_2545 (v820[11:0], v220[8:0], v2545[12:0]); // 3.0
    wire [11:0] v2546; shift_adder #(11, 11, 1, 1, 12, 0, 0) op_2546 (v821[10:0], v822[10:0], v2546[11:0]); // 3.0
    wire [14:0] v2547; shift_adder #(13, 12, 1, 1, 15, 2, 0) op_2547 (v823[12:0], v824[11:0], v2547[14:0]); // 3.0
    wire [12:0] v2548; shift_adder #(12, 13, 1, 1, 13, 0, 0) op_2548 (v825[11:0], v826[12:0], v2548[12:0]); // 3.0
    wire [14:0] v2549; shift_adder #(14, 13, 1, 1, 15, 2, 0) op_2549 (v827[13:0], v828[12:0], v2549[14:0]); // 3.0
    wire [19:0] v2550; shift_adder #(8, 16, 1, 1, 20, -11, 0) op_2550 (v116[7:0], v778[15:0], v2550[19:0]); // 3.0
    wire [26:0] v2551; shift_adder #(8, 25, 1, 1, 27, -18, 1) op_2551 (v84[7:0], v829[24:0], v2551[26:0]); // 3.0
    wire [13:0] v2552; shift_adder #(11, 14, 1, 1, 14, -1, 0) op_2552 (v228[10:0], v830[13:0], v2552[13:0]); // 3.0
    wire [23:0] v2553; shift_adder #(8, 12, 1, 1, 24, 12, 0) op_2553 (v106[7:0], v831[11:0], v2553[23:0]); // 3.0
    wire [17:0] v2554; shift_adder #(11, 17, 1, 1, 18, -7, 0) op_2554 (v232[10:0], v832[16:0], v2554[17:0]); // 3.0
    wire [14:0] v2555; shift_adder #(8, 13, 1, 1, 15, 2, 0) op_2555 (v103[7:0], v833[12:0], v2555[14:0]); // 3.0
    wire [17:0] v2556; shift_adder #(14, 13, 1, 1, 18, -4, 0) op_2556 (v236[13:0], v834[12:0], v2556[17:0]); // 3.0
    wire [16:0] v2557; shift_adder #(12, 16, 1, 1, 17, -4, 0) op_2557 (v835[11:0], v836[15:0], v2557[16:0]); // 3.0
    wire [27:0] v2558; shift_adder #(13, 27, 1, 1, 28, -14, 0) op_2558 (v837[12:0], v838[26:0], v2558[27:0]); // 3.0
    wire [16:0] v2559; shift_adder #(12, 15, 1, 1, 17, 2, 1) op_2559 (v243[11:0], v839[14:0], v2559[16:0]); // 3.0
    wire [19:0] v2560; shift_adder #(15, 20, 1, 1, 20, -3, 0) op_2560 (v840[14:0], v841[19:0], v2560[19:0]); // 3.0
    wire [16:0] v2561; shift_adder #(12, 14, 1, 1, 17, 3, 1) op_2561 (v247[11:0], v842[13:0], v2561[16:0]); // 3.0
    wire [22:0] v2562; shift_adder #(12, 22, 1, 1, 23, -10, 0) op_2562 (v843[11:0], v844[21:0], v2562[22:0]); // 3.0
    wire [21:0] v2563; shift_adder #(11, 13, 1, 1, 22, 9, 1) op_2563 (v177[10:0], v845[12:0], v2563[21:0]); // 3.0
    wire [15:0] v2564; shift_adder #(11, 10, 1, 1, 16, -5, 0) op_2564 (v846[10:0], v252[9:0], v2564[15:0]); // 3.0
    wire [17:0] v2565; shift_adder #(17, 12, 1, 1, 18, 5, 0) op_2565 (v847[16:0], v848[11:0], v2565[17:0]); // 3.0
    wire [15:0] v2566; shift_adder #(11, 16, 1, 1, 16, -4, 0) op_2566 (v134[10:0], v849[15:0], v2566[15:0]); // 3.0
    wire [30:0] v2567; shift_adder #(29, 23, 1, 1, 31, 7, 0) op_2567 (v850[28:0], v851[22:0], v2567[30:0]); // 3.0
    wire [28:0] v2568; shift_adder #(17, 19, 1, 1, 29, -12, 0) op_2568 (v852[16:0], v805[18:0], v2568[28:0]); // 3.0
    wire [17:0] v2569; shift_adder #(18, 12, 1, 1, 18, 4, 0) op_2569 (v853[17:0], v854[11:0], v2569[17:0]); // 3.0
    wire [17:0] v2570; shift_adder #(11, 18, 1, 1, 18, -6, 0) op_2570 (v855[10:0], v856[17:0], v2570[17:0]); // 3.0
    wire [33:0] v2571; shift_adder #(12, 33, 1, 1, 34, -21, 0) op_2571 (v857[11:0], v858[32:0], v2571[33:0]); // 3.0
    wire [12:0] v2572; shift_adder #(13, 10, 1, 1, 13, 0, 0) op_2572 (v859[12:0], v263[9:0], v2572[12:0]); // 3.0
    wire [15:0] v2573; shift_adder #(13, 13, 1, 1, 16, -3, 0) op_2573 (v860[12:0], v861[12:0], v2573[15:0]); // 3.0
    wire [13:0] v2574; shift_adder #(11, 12, 1, 1, 14, -3, 0) op_2574 (v193[10:0], v862[11:0], v2574[13:0]); // 3.0
    wire [12:0] v2575; shift_adder #(8, 12, 1, 1, 13, -4, 1) op_2575 (v72[7:0], v863[11:0], v2575[12:0]); // 3.0
    wire [30:0] v2576; shift_adder #(11, 24, 1, 1, 31, 7, 0) op_2576 (v268[10:0], v864[23:0], v2576[30:0]); // 3.0
    wire [18:0] v2577; shift_adder #(18, 15, 1, 1, 19, 3, 0) op_2577 (v865[17:0], v866[14:0], v2577[18:0]); // 3.0
    wire [14:0] v2578; shift_adder #(12, 14, 1, 1, 15, -2, 0) op_2578 (v867[11:0], v271[13:0], v2578[14:0]); // 3.0
    wire [16:0] v2579; shift_adder #(17, 11, 1, 1, 17, 3, 0) op_2579 (v869[16:0], v870[10:0], v2579[16:0]); // 3.0
    wire [17:0] v2580; shift_adder #(14, 18, 1, 1, 18, -2, 0) op_2580 (v871[13:0], v872[17:0], v2580[17:0]); // 3.0
    wire [17:0] v2581; shift_adder #(12, 18, 1, 1, 18, -3, 1) op_2581 (v873[11:0], v874[17:0], v2581[17:0]); // 3.0
    wire [17:0] v2582; shift_adder #(17, 17, 1, 1, 18, 1, 0) op_2582 (v875[16:0], v876[16:0], v2582[17:0]); // 3.0
    wire [14:0] v2583; shift_adder #(13, 14, 1, 1, 15, -1, 0) op_2583 (v877[12:0], v878[13:0], v2583[14:0]); // 3.0
    wire [18:0] v2584; shift_adder #(12, 13, 1, 1, 19, -7, 1) op_2584 (v285[11:0], v880[12:0], v2584[18:0]); // 3.0
    wire [18:0] v2585; shift_adder #(18, 17, 1, 1, 19, 2, 1) op_2585 (v286[17:0], v881[16:0], v2585[18:0]); // 3.0
    wire [13:0] v2586; shift_adder #(12, 13, 1, 1, 14, -2, 1) op_2586 (v288[11:0], v882[12:0], v2586[13:0]); // 3.0
    wire [21:0] v2587; shift_adder #(13, 10, 1, 1, 22, -9, 0) op_2587 (v883[12:0], v291[9:0], v2587[21:0]); // 3.0
    wire [12:0] v2588; shift_adder #(13, 11, 1, 1, 13, 0, 0) op_2588 (v884[12:0], v885[10:0], v2588[12:0]); // 3.0
    wire [17:0] v2589; shift_adder #(8, 15, 1, 1, 18, 3, 0) op_2589 (v127[7:0], v886[14:0], v2589[17:0]); // 3.0
    wire [19:0] v2590; shift_adder #(17, 15, 1, 1, 20, 5, 0) op_2590 (v887[16:0], v295[14:0], v2590[19:0]); // 3.0
    wire [16:0] v2591; shift_adder #(13, 17, 1, 1, 17, -2, 0) op_2591 (v888[12:0], v889[16:0], v2591[16:0]); // 3.0
    wire [20:0] v2592; shift_adder #(11, 17, 1, 1, 21, 4, 1) op_2592 (v178[10:0], v890[16:0], v2592[20:0]); // 3.0
    wire [14:0] v2593; shift_adder #(11, 13, 1, 1, 15, 2, 1) op_2593 (v181[10:0], v803[12:0], v2593[14:0]); // 3.0
    wire [14:0] v2594; shift_adder #(13, 13, 1, 1, 15, 2, 0) op_2594 (v891[12:0], v892[12:0], v2594[14:0]); // 3.0
    wire [15:0] v2595; shift_adder #(15, 15, 1, 1, 16, 0, 0) op_2595 (v893[14:0], v894[14:0], v2595[15:0]); // 3.0
    wire [19:0] v2596; shift_adder #(11, 17, 1, 1, 20, -9, 0) op_2596 (v228[10:0], v895[16:0], v2596[19:0]); // 3.0
    wire [17:0] v2597; shift_adder #(12, 17, 1, 1, 18, -4, 0) op_2597 (v896[11:0], v897[16:0], v2597[17:0]); // 3.0
    wire [14:0] v2598; shift_adder #(13, 14, 1, 1, 15, 0, 0) op_2598 (v898[12:0], v899[13:0], v2598[14:0]); // 3.0
    wire [17:0] v2599; shift_adder #(11, 13, 1, 1, 18, 5, 0) op_2599 (v245[10:0], v900[12:0], v2599[17:0]); // 3.0
    wire [16:0] v2600; shift_adder #(16, 15, 1, 1, 17, -1, 0) op_2600 (v901[15:0], v902[14:0], v2600[16:0]); // 3.0
    wire [19:0] v2601; shift_adder #(19, 15, 1, 1, 20, 4, 0) op_2601 (v903[18:0], v904[14:0], v2601[19:0]); // 3.0
    wire [19:0] v2602; shift_adder #(13, 15, 1, 1, 20, 5, 1) op_2602 (v833[12:0], v905[14:0], v2602[19:0]); // 3.0
    wire [26:0] v2603; shift_adder #(22, 21, 1, 1, 27, 6, 0) op_2603 (v906[21:0], v907[20:0], v2603[26:0]); // 3.0
    wire [21:0] v2604; shift_adder #(8, 22, 1, 1, 22, -2, 0) op_2604 (v85[7:0], v908[21:0], v2604[21:0]); // 3.0
    wire [21:0] v2605; shift_adder #(8, 22, 1, 1, 22, -7, 1) op_2605 (v97[7:0], v909[21:0], v2605[21:0]); // 3.0
    wire [19:0] v2606; shift_adder #(19, 19, 1, 1, 20, 0, 0) op_2606 (v910[18:0], v911[18:0], v2606[19:0]); // 3.0
    wire [27:0] v2607; shift_adder #(27, 15, 1, 1, 28, 13, 0) op_2607 (v912[26:0], v913[14:0], v2607[27:0]); // 3.0
    wire [16:0] v2608; shift_adder #(15, 13, 1, 1, 17, 4, 0) op_2608 (v914[14:0], v915[12:0], v2608[16:0]); // 3.0
    wire [34:0] v2609; shift_adder #(15, 25, 1, 1, 35, 10, 0) op_2609 (v313[14:0], v916[24:0], v2609[34:0]); // 3.0
    wire [21:0] v2610; shift_adder #(17, 22, 1, 1, 22, -4, 0) op_2610 (v917[16:0], v918[21:0], v2610[21:0]); // 3.0
    wire [17:0] v2611; shift_adder #(8, 12, 1, 1, 18, 6, 0) op_2611 (v114[7:0], v919[11:0], v2611[17:0]); // 3.0
    wire [12:0] v2612; shift_adder #(8, 13, 1, 1, 13, 0, 1) op_2612 (v75[7:0], v860[12:0], v2612[12:0]); // 3.0
    wire [17:0] v2613; shift_adder #(13, 17, 1, 1, 18, -5, 0) op_2613 (v920[12:0], v921[16:0], v2613[17:0]); // 3.0
    wire [15:0] v2614; shift_adder #(11, 13, 1, 1, 16, -5, 0) op_2614 (v229[10:0], v837[12:0], v2614[15:0]); // 3.0
    wire [16:0] v2615; shift_adder #(15, 13, 1, 1, 17, -2, 1) op_2615 (v922[14:0], v923[12:0], v2615[16:0]); // 3.0
    wire [22:0] v2616; shift_adder #(11, 12, 1, 1, 23, -12, 0) op_2616 (v319[10:0], v924[11:0], v2616[22:0]); // 3.0
    wire [24:0] v2617; shift_adder #(17, 20, 1, 1, 25, 5, 1) op_2617 (v876[16:0], v925[19:0], v2617[24:0]); // 3.0
    wire [18:0] v2618; shift_adder #(18, 16, 1, 1, 19, 2, 0) op_2618 (v926[17:0], v927[15:0], v2618[18:0]); // 3.0
    wire [14:0] v2619; shift_adder #(14, 12, 1, 1, 15, 3, 0) op_2619 (v928[13:0], v929[11:0], v2619[14:0]); // 3.0
    wire [26:0] v2620; shift_adder #(8, 27, 1, 1, 27, -14, 1) op_2620 (v81[7:0], v930[26:0], v2620[26:0]); // 3.0
    wire [21:0] v2621; shift_adder #(8, 19, 1, 1, 22, -13, 1) op_2621 (v77[7:0], v931[18:0], v2621[21:0]); // 3.0
    wire [14:0] v2622; shift_adder #(8, 13, 1, 1, 15, -6, 1) op_2622 (v122[7:0], v932[12:0], v2622[14:0]); // 3.0
    wire [26:0] v2623; shift_adder #(14, 27, 1, 1, 27, -6, 0) op_2623 (v830[13:0], v933[26:0], v2623[26:0]); // 3.0
    wire [25:0] v2624; shift_adder #(12, 12, 1, 1, 26, -14, 0) op_2624 (v934[11:0], v935[11:0], v2624[25:0]); // 3.0
    wire [14:0] v2625; shift_adder #(11, 12, 1, 1, 15, -4, 0) op_2625 (v147[10:0], v936[11:0], v2625[14:0]); // 3.0
    wire [17:0] v2626; shift_adder #(14, 18, 1, 1, 18, -3, 0) op_2626 (v937[13:0], v938[17:0], v2626[17:0]); // 3.0
    wire [18:0] v2627; shift_adder #(18, 18, 1, 1, 19, -1, 0) op_2627 (v939[17:0], v940[17:0], v2627[18:0]); // 3.0
    wire [20:0] v2628; shift_adder #(11, 11, 1, 1, 21, -10, 1) op_2628 (v941[10:0], v330[10:0], v2628[20:0]); // 3.0
    wire [21:0] v2629; shift_adder #(12, 21, 1, 1, 22, -10, 0) op_2629 (v942[11:0], v943[20:0], v2629[21:0]); // 3.0
    wire [20:0] v2630; shift_adder #(19, 15, 1, 1, 21, -2, 1) op_2630 (v944[18:0], v945[14:0], v2630[20:0]); // 3.0
    wire [33:0] v2631; shift_adder #(16, 32, 1, 1, 34, -17, 0) op_2631 (v946[15:0], v947[31:0], v2631[33:0]); // 3.0
    wire [25:0] v2632; shift_adder #(12, 13, 1, 1, 26, -14, 0) op_2632 (v333[11:0], v948[12:0], v2632[25:0]); // 3.0
    wire [17:0] v2633; shift_adder #(18, 14, 1, 1, 18, 3, 0) op_2633 (v949[17:0], v950[13:0], v2633[17:0]); // 3.0
    wire [25:0] v2634; shift_adder #(13, 21, 1, 1, 26, 5, 1) op_2634 (v149[12:0], v951[20:0], v2634[25:0]); // 3.0
    wire [17:0] v2635; shift_adder #(17, 13, 1, 1, 18, 5, 0) op_2635 (v952[16:0], v953[12:0], v2635[17:0]); // 3.0
    wire [34:0] v2636; shift_adder #(11, 34, 1, 1, 35, -23, 0) op_2636 (v954[10:0], v955[33:0], v2636[34:0]); // 3.0
    wire [15:0] v2637; shift_adder #(12, 12, 1, 1, 16, -3, 0) op_2637 (v956[11:0], v957[11:0], v2637[15:0]); // 3.0
    wire [13:0] v2638; shift_adder #(8, 14, 1, 1, 14, -2, 1) op_2638 (v92[7:0], v958[13:0], v2638[13:0]); // 3.0
    wire [15:0] v2639; shift_adder #(16, 14, 1, 1, 16, 0, 0) op_2639 (v959[15:0], v960[13:0], v2639[15:0]); // 3.0
    wire [17:0] v2640; shift_adder #(8, 11, 1, 1, 18, -9, 0) op_2640 (v122[7:0], v961[10:0], v2640[17:0]); // 3.0
    wire [16:0] v2641; shift_adder #(13, 11, 1, 1, 17, -4, 1) op_2641 (v346[12:0], v962[10:0], v2641[16:0]); // 3.0
    wire [16:0] v2642; shift_adder #(17, 14, 1, 1, 17, 1, 0) op_2642 (v963[16:0], v964[13:0], v2642[16:0]); // 3.0
    wire [16:0] v2643; shift_adder #(11, 12, 1, 1, 17, -6, 1) op_2643 (v134[10:0], v965[11:0], v2643[16:0]); // 3.0
    wire [17:0] v2644; shift_adder #(13, 17, 1, 1, 18, -4, 0) op_2644 (v790[12:0], v966[16:0], v2644[17:0]); // 3.0
    wire [17:0] v2645; shift_adder #(13, 17, 1, 1, 18, -5, 0) op_2645 (v882[12:0], v967[16:0], v2645[17:0]); // 3.0
    wire [20:0] v2646; shift_adder #(9, 18, 1, 1, 21, -11, 0) op_2646 (v351[8:0], v874[17:0], v2646[20:0]); // 3.0
    wire [19:0] v2647; shift_adder #(11, 18, 1, 1, 20, 2, 0) op_2647 (v329[10:0], v968[17:0], v2647[19:0]); // 3.0
    wire [20:0] v2648; shift_adder #(8, 15, 1, 1, 21, -12, 0) op_2648 (v70[7:0], v969[14:0], v2648[20:0]); // 3.0
    wire [15:0] v2649; shift_adder #(16, 12, 1, 1, 16, 3, 0) op_2649 (v970[15:0], v971[11:0], v2649[15:0]); // 3.0
    wire [17:0] v2650; shift_adder #(17, 12, 1, 1, 18, 5, 0) op_2650 (v972[16:0], v973[11:0], v2650[17:0]); // 3.0
    wire [13:0] v2651; shift_adder #(13, 14, 1, 1, 14, 0, 0) op_2651 (v974[12:0], v975[13:0], v2651[13:0]); // 3.0
    wire [14:0] v2652; shift_adder #(13, 14, 1, 1, 15, 0, 0) op_2652 (v900[12:0], v976[13:0], v2652[14:0]); // 3.0
    wire [18:0] v2653; shift_adder #(11, 19, 1, 1, 19, -2, 0) op_2653 (v187[10:0], v944[18:0], v2653[18:0]); // 3.0
    wire [18:0] v2654; shift_adder #(18, 13, 1, 1, 19, 5, 0) op_2654 (v977[17:0], v978[12:0], v2654[18:0]); // 3.0
    wire [27:0] v2655; shift_adder #(26, 23, 1, 1, 28, 4, 0) op_2655 (v979[25:0], v980[22:0], v2655[27:0]); // 3.0
    wire [17:0] v2656; shift_adder #(12, 17, 1, 1, 18, -6, 0) op_2656 (v981[11:0], v982[16:0], v2656[17:0]); // 3.0
    wire [16:0] v2657; shift_adder #(11, 17, 1, 1, 17, -5, 1) op_2657 (v284[10:0], v852[16:0], v2657[16:0]); // 3.0
    wire [18:0] v2658; shift_adder #(8, 13, 1, 1, 19, -10, 0) op_2658 (v85[7:0], v880[12:0], v2658[18:0]); // 3.0
    wire [37:0] v2659; shift_adder #(13, 14, 1, 1, 38, 24, 1) op_2659 (v983[12:0], v356[13:0], v2659[37:0]); // 3.0
    wire [30:0] v2660; shift_adder #(30, 13, 1, 1, 31, 17, 0) op_2660 (v984[29:0], v985[12:0], v2660[30:0]); // 3.0
    wire [15:0] v2661; shift_adder #(14, 11, 1, 1, 16, 4, 0) op_2661 (v986[13:0], v987[10:0], v2661[15:0]); // 3.0
    wire [18:0] v2662; shift_adder #(18, 12, 1, 1, 19, 6, 0) op_2662 (v989[17:0], v867[11:0], v2662[18:0]); // 3.0
    wire [13:0] v2663; shift_adder #(12, 12, 1, 1, 14, -1, 0) op_2663 (v990[11:0], v991[11:0], v2663[13:0]); // 3.0
    wire [13:0] v2664; shift_adder #(11, 13, 1, 1, 14, 1, 1) op_2664 (v251[10:0], v833[12:0], v2664[13:0]); // 3.0
    wire [15:0] v2665; shift_adder #(14, 15, 1, 1, 16, -1, 0) op_2665 (v992[13:0], v993[14:0], v2665[15:0]); // 3.0
    wire [22:0] v2666; shift_adder #(23, 17, 1, 1, 23, 5, 1) op_2666 (v258[22:0], v773[16:0], v2666[22:0]); // 3.0
    wire [22:0] v2667; shift_adder #(17, 21, 1, 1, 23, -6, 0) op_2667 (v921[16:0], v994[20:0], v2667[22:0]); // 3.0
    wire [18:0] v2668; shift_adder #(13, 13, 1, 1, 19, -6, 1) op_2668 (v995[12:0], v996[12:0], v2668[18:0]); // 3.0
    wire [22:0] v2669; shift_adder #(14, 21, 1, 1, 23, -8, 0) op_2669 (v997[13:0], v998[20:0], v2669[22:0]); // 3.0
    wire [18:0] v2670; shift_adder #(9, 12, 1, 1, 19, 7, 1) op_2670 (v360[8:0], v999[11:0], v2670[18:0]); // 3.0
    wire [18:0] v2671; shift_adder #(11, 12, 1, 1, 19, 7, 1) op_2671 (v268[10:0], v1000[11:0], v2671[18:0]); // 3.0
    wire [13:0] v2672; shift_adder #(13, 14, 1, 1, 14, 0, 0) op_2672 (v1001[12:0], v1002[13:0], v2672[13:0]); // 3.0
    wire [22:0] v2673; shift_adder #(22, 12, 1, 1, 23, 10, 0) op_2673 (v1003[21:0], v934[11:0], v2673[22:0]); // 3.0
    wire [12:0] v2674; shift_adder #(11, 12, 1, 1, 13, 1, 0) op_2674 (v367[10:0], v1004[11:0], v2674[12:0]); // 3.0
    wire [24:0] v2675; shift_adder #(16, 18, 1, 1, 25, -9, 1) op_2675 (v927[15:0], v1005[17:0], v2675[24:0]); // 3.0
    wire [16:0] v2676; shift_adder #(9, 15, 1, 1, 17, 2, 0) op_2676 (v369[8:0], v1006[14:0], v2676[16:0]); // 3.0
    wire [22:0] v2677; shift_adder #(14, 22, 1, 1, 23, -8, 0) op_2677 (v1007[13:0], v1008[21:0], v2677[22:0]); // 3.0
    wire [18:0] v2678; shift_adder #(12, 19, 1, 1, 19, -1, 1) op_2678 (v372[11:0], v1009[18:0], v2678[18:0]); // 3.0
    wire [25:0] v2679; shift_adder #(15, 26, 1, 1, 26, 0, 1) op_2679 (v1010[14:0], v373[25:0], v2679[25:0]); // 3.0
    wire [15:0] v2680; shift_adder #(15, 15, 1, 1, 16, -1, 0) op_2680 (v1011[14:0], v1012[14:0], v2680[15:0]); // 3.0
    wire [29:0] v2681; shift_adder #(14, 14, 1, 1, 30, -16, 0) op_2681 (v1013[13:0], v1014[13:0], v2681[29:0]); // 3.0
    wire [21:0] v2682; shift_adder #(13, 19, 1, 1, 22, 3, 1) op_2682 (v845[12:0], v376[18:0], v2682[21:0]); // 3.0
    wire [22:0] v2683; shift_adder #(15, 17, 1, 1, 23, 6, 1) op_2683 (v1015[14:0], v1016[16:0], v2683[22:0]); // 3.0
    wire [24:0] v2684; shift_adder #(25, 13, 1, 1, 25, 10, 0) op_2684 (v1017[24:0], v1018[12:0], v2684[24:0]); // 3.0
    wire [15:0] v2685; shift_adder #(11, 15, 1, 1, 16, -4, 0) op_2685 (v148[10:0], v1019[14:0], v2685[15:0]); // 3.0
    wire [16:0] v2686; shift_adder #(11, 16, 1, 1, 17, 1, 1) op_2686 (v379[10:0], v1020[15:0], v2686[16:0]); // 3.0
    wire [33:0] v2687; shift_adder #(13, 11, 1, 1, 34, -21, 1) op_2687 (v1021[12:0], v885[10:0], v2687[33:0]); // 3.0
    wire [30:0] v2688; shift_adder #(28, 17, 1, 1, 31, 14, 0) op_2688 (v1022[27:0], v1023[16:0], v2688[30:0]); // 3.0
    wire [13:0] v2689; shift_adder #(13, 12, 1, 1, 14, -1, 0) op_2689 (v1024[12:0], v1025[11:0], v2689[13:0]); // 3.0
    wire [17:0] v2690; shift_adder #(11, 13, 1, 1, 18, 5, 0) op_2690 (v131[10:0], v1026[12:0], v2690[17:0]); // 3.0
    wire [17:0] v2691; shift_adder #(15, 16, 1, 1, 18, 2, 0) op_2691 (v1027[14:0], v1028[15:0], v2691[17:0]); // 3.0
    wire [13:0] v2692; shift_adder #(13, 13, 1, 1, 14, -1, 0) op_2692 (v1029[12:0], v1030[12:0], v2692[13:0]); // 3.0
    wire [21:0] v2693; shift_adder #(12, 12, 1, 1, 22, 10, 0) op_2693 (v383[11:0], v1031[11:0], v2693[21:0]); // 3.0
    wire [14:0] v2694; shift_adder #(11, 13, 1, 1, 15, -4, 1) op_2694 (v328[10:0], v995[12:0], v2694[14:0]); // 3.0
    wire [19:0] v2695; shift_adder #(18, 16, 1, 1, 20, 4, 0) op_2695 (v1032[17:0], v1033[15:0], v2695[19:0]); // 3.0
    wire [16:0] v2696; shift_adder #(13, 12, 1, 1, 17, -4, 1) op_2696 (v1034[12:0], v1035[11:0], v2696[16:0]); // 3.0
    wire [18:0] v2697; shift_adder #(19, 17, 1, 1, 19, 1, 0) op_2697 (v1036[18:0], v1037[16:0], v2697[18:0]); // 3.0
    wire [21:0] v2698; shift_adder #(11, 15, 1, 1, 22, 7, 1) op_2698 (v289[10:0], v1038[14:0], v2698[21:0]); // 3.0
    wire [20:0] v2699; shift_adder #(14, 21, 1, 1, 21, -6, 0) op_2699 (v1039[13:0], v1040[20:0], v2699[20:0]); // 3.0
    wire [25:0] v2700; shift_adder #(13, 13, 1, 1, 26, 13, 0) op_2700 (v883[12:0], v1041[12:0], v2700[25:0]); // 3.0
    wire [25:0] v2701; shift_adder #(26, 13, 1, 1, 26, 10, 0) op_2701 (v1042[25:0], v948[12:0], v2701[25:0]); // 3.0
    wire [24:0] v2702; shift_adder #(12, 24, 1, 1, 25, -13, 1) op_2702 (v1043[11:0], v1044[23:0], v2702[24:0]); // 3.0
    wire [13:0] v2703; shift_adder #(13, 13, 1, 1, 14, 0, 0) op_2703 (v1021[12:0], v1029[12:0], v2703[13:0]); // 3.0
    wire [14:0] v2704; shift_adder #(8, 14, 1, 1, 15, 1, 0) op_2704 (v116[7:0], v1045[13:0], v2704[14:0]); // 3.0
    wire [14:0] v2705; shift_adder #(13, 12, 1, 1, 15, 3, 0) op_2705 (v1046[12:0], v1047[11:0], v2705[14:0]); // 3.0
    wire [25:0] v2706; shift_adder #(11, 26, 1, 1, 26, -13, 0) op_2706 (v1049[10:0], v1050[25:0], v2706[25:0]); // 3.0
    wire [33:0] v2707; shift_adder #(33, 15, 1, 1, 34, 19, 0) op_2707 (v1051[32:0], v1052[14:0], v2707[33:0]); // 3.0
    wire [15:0] v2708; shift_adder #(15, 11, 1, 1, 16, 4, 0) op_2708 (v1053[14:0], v1054[10:0], v2708[15:0]); // 3.0
    wire [14:0] v2709; shift_adder #(11, 12, 1, 1, 15, 3, 0) op_2709 (v393[10:0], v879[11:0], v2709[14:0]); // 3.0
    wire [14:0] v2710; shift_adder #(8, 15, 1, 1, 15, -2, 0) op_2710 (v79[7:0], v1055[14:0], v2710[14:0]); // 3.0
    wire [15:0] v2711; shift_adder #(12, 14, 1, 1, 16, -3, 0) op_2711 (v1056[11:0], v1057[13:0], v2711[15:0]); // 3.0
    wire [31:0] v2712; shift_adder #(9, 24, 1, 1, 32, -22, 0) op_2712 (v395[8:0], v1058[23:0], v2712[31:0]); // 3.0
    wire [32:0] v2713; shift_adder #(19, 33, 1, 1, 33, -13, 0) op_2713 (v1059[18:0], v1060[32:0], v2713[32:0]); // 3.0
    wire [22:0] v2714; shift_adder #(8, 22, 1, 1, 23, -13, 0) op_2714 (v95[7:0], v1061[21:0], v2714[22:0]); // 3.0
    wire [24:0] v2715; shift_adder #(13, 21, 1, 1, 25, 4, 0) op_2715 (v189[12:0], v1062[20:0], v2715[24:0]); // 3.0
    wire [20:0] v2716; shift_adder #(17, 16, 1, 1, 21, 5, 0) op_2716 (v1063[16:0], v1064[15:0], v2716[20:0]); // 3.0
    wire [35:0] v2717; shift_adder #(35, 15, 1, 1, 36, 20, 0) op_2717 (v1065[34:0], v1066[14:0], v2717[35:0]); // 3.0
    wire [22:0] v2718; shift_adder #(22, 12, 1, 1, 23, 10, 0) op_2718 (v1067[21:0], v1068[11:0], v2718[22:0]); // 3.0
    wire [13:0] v2719; shift_adder #(8, 12, 1, 1, 14, -5, 1) op_2719 (v66[7:0], v1069[11:0], v2719[13:0]); // 3.0
    wire [15:0] v2720; shift_adder #(13, 15, 1, 1, 16, -2, 0) op_2720 (v1070[12:0], v1071[14:0], v2720[15:0]); // 3.0
    wire [14:0] v2721; shift_adder #(12, 13, 1, 1, 15, -3, 1) op_2721 (v397[11:0], v915[12:0], v2721[14:0]); // 3.0
    wire [18:0] v2722; shift_adder #(14, 18, 1, 1, 19, -4, 0) op_2722 (v1072[13:0], v1073[17:0], v2722[18:0]); // 3.0
    wire [19:0] v2723; shift_adder #(13, 20, 1, 1, 20, -2, 1) op_2723 (v1074[12:0], v1075[19:0], v2723[19:0]); // 3.0
    wire [26:0] v2724; shift_adder #(12, 26, 1, 1, 27, -15, 0) op_2724 (v404[11:0], v1076[25:0], v2724[26:0]); // 3.0
    wire [12:0] v2725; shift_adder #(12, 12, 1, 1, 13, 0, 0) op_2725 (v862[11:0], v1077[11:0], v2725[12:0]); // 3.0
    wire [17:0] v2726; shift_adder #(12, 13, 1, 1, 18, -6, 1) op_2726 (v321[11:0], v1078[12:0], v2726[17:0]); // 3.0
    wire [17:0] v2727; shift_adder #(13, 16, 1, 1, 18, -5, 0) op_2727 (v1079[12:0], v901[15:0], v2727[17:0]); // 3.0
    wire [12:0] v2728; shift_adder #(12, 11, 1, 1, 13, 0, 0) op_2728 (v1080[11:0], v1081[10:0], v2728[12:0]); // 3.0
    wire [13:0] v2729; shift_adder #(12, 13, 1, 1, 14, -2, 0) op_2729 (v1082[11:0], v406[12:0], v2729[13:0]); // 3.0
    wire [15:0] v2730; shift_adder #(13, 15, 1, 1, 16, -3, 0) op_2730 (v1083[12:0], v1084[14:0], v2730[15:0]); // 3.0
    wire [14:0] v2731; shift_adder #(14, 14, 1, 1, 15, 1, 0) op_2731 (v830[13:0], v1085[13:0], v2731[14:0]); // 3.0
    wire [13:0] v2732; shift_adder #(13, 13, 1, 1, 14, -1, 0) op_2732 (v793[12:0], v1086[12:0], v2732[13:0]); // 3.0
    wire [11:0] v2733; shift_adder #(8, 11, 1, 1, 12, -1, 1) op_2733 (v77[7:0], v846[10:0], v2733[11:0]); // 3.0
    wire [26:0] v2734; shift_adder #(24, 16, 1, 1, 27, 11, 0) op_2734 (v1087[23:0], v1088[15:0], v2734[26:0]); // 3.0
    wire [20:0] v2735; shift_adder #(13, 13, 1, 1, 21, 8, 1) op_2735 (v932[12:0], v1079[12:0], v2735[20:0]); // 3.0
    wire [26:0] v2736; shift_adder #(8, 16, 1, 1, 27, 11, 1) op_2736 (v90[7:0], v1089[15:0], v2736[26:0]); // 3.0
    wire [20:0] v2737; shift_adder #(21, 16, 1, 1, 21, 2, 0) op_2737 (v1090[20:0], v1091[15:0], v2737[20:0]); // 3.0
    wire [29:0] v2738; shift_adder #(25, 30, 1, 1, 30, -4, 0) op_2738 (v1092[24:0], v1093[29:0], v2738[29:0]); // 3.0
    wire [19:0] v2739; shift_adder #(16, 18, 1, 1, 20, -4, 0) op_2739 (v901[15:0], v1094[17:0], v2739[19:0]); // 3.0
    wire [24:0] v2740; shift_adder #(19, 25, 1, 1, 25, -5, 0) op_2740 (v931[18:0], v1095[24:0], v2740[24:0]); // 3.0
    wire [30:0] v2741; shift_adder #(8, 27, 1, 1, 31, -22, 0) op_2741 (v107[7:0], v838[26:0], v2741[30:0]); // 3.0
    wire [31:0] v2742; shift_adder #(26, 18, 1, 1, 32, -6, 1) op_2742 (v373[25:0], v1096[17:0], v2742[31:0]); // 3.0
    wire [27:0] v2743; shift_adder #(11, 13, 1, 1, 28, 15, 0) op_2743 (v209[10:0], v1097[12:0], v2743[27:0]); // 3.0
    wire [17:0] v2744; shift_adder #(16, 18, 1, 1, 18, 0, 0) op_2744 (v1098[15:0], v1099[17:0], v2744[17:0]); // 3.0
    wire [12:0] v2745; shift_adder #(11, 12, 1, 1, 13, -1, 1) op_2745 (v136[10:0], v1100[11:0], v2745[12:0]); // 3.0
    wire [20:0] v2746; shift_adder #(12, 20, 1, 1, 21, -9, 0) op_2746 (v174[11:0], v1101[19:0], v2746[20:0]); // 3.0
    wire [14:0] v2747; shift_adder #(8, 12, 1, 1, 15, 3, 0) op_2747 (v88[7:0], v1102[11:0], v2747[14:0]); // 3.0
    wire [13:0] v2748; shift_adder #(12, 14, 1, 1, 14, 0, 0) op_2748 (v1103[11:0], v1104[13:0], v2748[13:0]); // 3.0
    wire [17:0] v2749; shift_adder #(11, 18, 1, 1, 18, -5, 0) op_2749 (v375[10:0], v865[17:0], v2749[17:0]); // 3.0
    wire [14:0] v2750; shift_adder #(12, 14, 1, 1, 15, -1, 0) op_2750 (v1105[11:0], v992[13:0], v2750[14:0]); // 3.0
    wire [20:0] v2751; shift_adder #(13, 16, 1, 1, 21, -8, 1) op_2751 (v416[12:0], v1106[15:0], v2751[20:0]); // 3.0
    wire [17:0] v2752; shift_adder #(15, 15, 1, 1, 18, 3, 0) op_2752 (v1107[14:0], v1108[14:0], v2752[17:0]); // 3.0
    wire [15:0] v2753; shift_adder #(15, 12, 1, 1, 16, 3, 0) op_2753 (v1109[14:0], v1068[11:0], v2753[15:0]); // 3.0
    wire [34:0] v2754; shift_adder #(34, 14, 1, 1, 35, 21, 0) op_2754 (v1110[33:0], v1111[13:0], v2754[34:0]); // 3.0
    wire [19:0] v2755; shift_adder #(14, 19, 1, 1, 20, -4, 0) op_2755 (v1112[13:0], v1113[18:0], v2755[19:0]); // 3.0
    wire [25:0] v2756; shift_adder #(11, 16, 1, 1, 26, 10, 0) op_2756 (v418[10:0], v1114[15:0], v2756[25:0]); // 3.0
    wire [14:0] v2757; shift_adder #(11, 14, 1, 1, 15, 1, 0) op_2757 (v1115[10:0], v1116[13:0], v2757[14:0]); // 3.0
    wire [14:0] v2758; shift_adder #(8, 14, 1, 1, 15, -6, 0) op_2758 (v68[7:0], v1117[13:0], v2758[14:0]); // 3.0
    wire [19:0] v2759; shift_adder #(17, 15, 1, 1, 20, -3, 1) op_2759 (v1118[16:0], v1119[14:0], v2759[19:0]); // 3.0
    wire [15:0] v2760; shift_adder #(15, 12, 1, 1, 16, 3, 0) op_2760 (v1120[14:0], v1121[11:0], v2760[15:0]); // 3.0
    wire [17:0] v2761; shift_adder #(11, 11, 1, 1, 18, 7, 0) op_2761 (v147[10:0], v1122[10:0], v2761[17:0]); // 3.0
    wire [13:0] v2762; shift_adder #(12, 13, 1, 1, 14, -1, 0) op_2762 (v285[11:0], v883[12:0], v2762[13:0]); // 3.0
    wire [14:0] v2763; shift_adder #(13, 15, 1, 1, 15, 0, 0) op_2763 (v1123[12:0], v1124[14:0], v2763[14:0]); // 3.0
    wire [17:0] v2764; shift_adder #(16, 13, 1, 1, 18, -2, 1) op_2764 (v426[15:0], v795[12:0], v2764[17:0]); // 3.0
    wire [14:0] v2765; shift_adder #(11, 12, 1, 1, 15, 2, 0) op_2765 (v147[10:0], v1125[11:0], v2765[14:0]); // 3.0
    wire [16:0] v2766; shift_adder #(14, 15, 1, 1, 17, 2, 0) op_2766 (v1126[13:0], v1127[14:0], v2766[16:0]); // 3.0
    wire [20:0] v2767; shift_adder #(8, 21, 1, 1, 21, -4, 1) op_2767 (v88[7:0], v1128[20:0], v2767[20:0]); // 3.0
    wire [16:0] v2768; shift_adder #(11, 13, 1, 1, 17, 4, 0) op_2768 (v203[10:0], v1030[12:0], v2768[16:0]); // 3.0
    wire [18:0] v2769; shift_adder #(15, 18, 1, 1, 19, -2, 0) op_2769 (v1129[14:0], v1130[17:0], v2769[18:0]); // 3.0
    wire [21:0] v2770; shift_adder #(19, 10, 1, 1, 22, -3, 0) op_2770 (v782[18:0], v263[9:0], v2770[21:0]); // 3.0
    wire [22:0] v2771; shift_adder #(23, 14, 1, 1, 23, 1, 0) op_2771 (v1131[22:0], v1132[13:0], v2771[22:0]); // 3.0
    wire [23:0] v2772; shift_adder #(22, 13, 1, 1, 24, 10, 0) op_2772 (v1133[21:0], v1134[12:0], v2772[23:0]); // 3.0
    wire [18:0] v2773; shift_adder #(11, 14, 1, 1, 19, 5, 0) op_2773 (v353[10:0], v1135[13:0], v2773[18:0]); // 3.0
    wire [18:0] v2774; shift_adder #(12, 13, 1, 1, 19, 6, 1) op_2774 (v1136[11:0], v923[12:0], v2774[18:0]); // 3.0
    wire [13:0] v2775; shift_adder #(11, 13, 1, 1, 14, -1, 0) op_2775 (v1137[10:0], v1138[12:0], v2775[13:0]); // 3.0
    wire [13:0] v2776; shift_adder #(11, 14, 1, 1, 14, 0, 1) op_2776 (v234[10:0], v1139[13:0], v2776[13:0]); // 3.0
    wire [30:0] v2777; shift_adder #(11, 31, 1, 1, 31, -9, 0) op_2777 (v141[10:0], v1140[30:0], v2777[30:0]); // 3.0
    wire [23:0] v2778; shift_adder #(23, 20, 1, 1, 24, 4, 1) op_2778 (v1141[22:0], v1142[19:0], v2778[23:0]); // 3.0
    wire [20:0] v2779; shift_adder #(19, 14, 1, 1, 21, 6, 0) op_2779 (v1143[18:0], v975[13:0], v2779[20:0]); // 3.0
    wire [23:0] v2780; shift_adder #(14, 23, 1, 1, 24, -9, 0) op_2780 (v1007[13:0], v788[22:0], v2780[23:0]); // 3.0
    wire [23:0] v2781; shift_adder #(21, 15, 1, 1, 24, -3, 0) op_2781 (v1144[20:0], v431[14:0], v2781[23:0]); // 3.0
    wire [30:0] v2782; shift_adder #(8, 31, 1, 1, 31, -14, 1) op_2782 (v89[7:0], v1145[30:0], v2782[30:0]); // 3.0
    wire [13:0] v2783; shift_adder #(11, 12, 1, 1, 14, -3, 0) op_2783 (v218[10:0], v1147[11:0], v2783[13:0]); // 3.0
    wire [24:0] v2784; shift_adder #(21, 24, 1, 1, 25, -3, 0) op_2784 (v1148[20:0], v1149[23:0], v2784[24:0]); // 3.0
    wire [23:0] v2785; shift_adder #(22, 18, 1, 1, 24, 6, 0) op_2785 (v1008[21:0], v1150[17:0], v2785[23:0]); // 3.0
    wire [18:0] v2786; shift_adder #(17, 16, 1, 1, 19, -2, 1) op_2786 (v1151[16:0], v1152[15:0], v2786[18:0]); // 3.0
    wire [15:0] v2787; shift_adder #(8, 12, 1, 1, 16, 4, 0) op_2787 (v87[7:0], v956[11:0], v2787[15:0]); // 3.0
    wire [13:0] v2788; shift_adder #(11, 12, 1, 1, 14, 1, 1) op_2788 (v319[10:0], v1153[11:0], v2788[13:0]); // 3.0
    wire [27:0] v2789; shift_adder #(8, 17, 1, 1, 28, 11, 1) op_2789 (v75[7:0], v1154[16:0], v2789[27:0]); // 3.0
    wire [16:0] v2790; shift_adder #(12, 16, 1, 1, 17, -4, 0) op_2790 (v1155[11:0], v1156[15:0], v2790[16:0]); // 3.0
    wire [18:0] v2791; shift_adder #(17, 15, 1, 1, 19, 3, 0) op_2791 (v1157[16:0], v1158[14:0], v2791[18:0]); // 3.0
    wire [36:0] v2792; shift_adder #(12, 14, 1, 1, 37, -25, 1) op_2792 (v862[11:0], v950[13:0], v2792[36:0]); // 3.0
    wire [13:0] v2793; shift_adder #(12, 12, 1, 1, 14, -1, 0) op_2793 (v1159[11:0], v1160[11:0], v2793[13:0]); // 3.0
    wire [14:0] v2794; shift_adder #(11, 13, 1, 1, 15, -4, 1) op_2794 (v1161[10:0], v272[12:0], v2794[14:0]); // 3.0
    wire [14:0] v2795; shift_adder #(11, 14, 1, 1, 15, 1, 1) op_2795 (v324[10:0], v1162[13:0], v2795[14:0]); // 3.0
    wire [14:0] v2796; shift_adder #(13, 13, 1, 1, 15, -2, 0) op_2796 (v1163[12:0], v1164[12:0], v2796[14:0]); // 3.0
    wire [18:0] v2797; shift_adder #(12, 14, 1, 1, 19, 5, 1) op_2797 (v411[11:0], v1165[13:0], v2797[18:0]); // 3.0
    wire [28:0] v2798; shift_adder #(11, 29, 1, 1, 29, -8, 1) op_2798 (v153[10:0], v1166[28:0], v2798[28:0]); // 3.0
    wire [25:0] v2799; shift_adder #(26, 21, 1, 1, 26, 4, 0) op_2799 (v1167[25:0], v1168[20:0], v2799[25:0]); // 3.0
    wire [31:0] v2800; shift_adder #(11, 16, 1, 1, 32, 16, 0) op_2800 (v241[10:0], v1169[15:0], v2800[31:0]); // 3.0
    wire [16:0] v2801; shift_adder #(11, 12, 1, 1, 17, 5, 0) op_2801 (v413[10:0], v1170[11:0], v2801[16:0]); // 3.0
    wire [18:0] v2802; shift_adder #(8, 12, 1, 1, 19, 7, 0) op_2802 (v85[7:0], v1171[11:0], v2802[18:0]); // 3.0
    wire [24:0] v2803; shift_adder #(17, 24, 1, 1, 25, -8, 0) op_2803 (v881[16:0], v1172[23:0], v2803[24:0]); // 3.0
    wire [16:0] v2804; shift_adder #(11, 15, 1, 1, 17, 2, 0) op_2804 (v228[10:0], v1173[14:0], v2804[16:0]); // 3.0
    wire [17:0] v2805; shift_adder #(11, 17, 1, 1, 18, -5, 0) op_2805 (v1174[10:0], v1175[16:0], v2805[17:0]); // 3.0
    wire [13:0] v2806; shift_adder #(12, 13, 1, 1, 14, -1, 0) op_2806 (v1176[11:0], v1177[12:0], v2806[13:0]); // 3.0
    wire [21:0] v2807; shift_adder #(12, 22, 1, 1, 22, -7, 0) op_2807 (v1178[11:0], v1179[21:0], v2807[21:0]); // 3.0
    wire [21:0] v2808; shift_adder #(13, 21, 1, 1, 22, -7, 0) op_2808 (v1180[12:0], v1181[20:0], v2808[21:0]); // 3.0
    wire [17:0] v2809; shift_adder #(12, 15, 1, 1, 18, -5, 0) op_2809 (v1182[11:0], v1183[14:0], v2809[17:0]); // 3.0
    wire [13:0] v2810; shift_adder #(13, 11, 1, 1, 14, 1, 0) op_2810 (v1184[12:0], v1185[10:0], v2810[13:0]); // 3.0
    wire [15:0] v2811; shift_adder #(15, 13, 1, 1, 16, 2, 0) op_2811 (v1186[14:0], v1187[12:0], v2811[15:0]); // 3.0
    wire [31:0] v2812; shift_adder #(8, 12, 1, 1, 32, -23, 0) op_2812 (v114[7:0], v1188[11:0], v2812[31:0]); // 3.0
    wire [23:0] v2813; shift_adder #(13, 10, 1, 1, 24, 14, 0) op_2813 (v1189[12:0], v446[9:0], v2813[23:0]); // 3.0
    wire [34:0] v2814; shift_adder #(12, 12, 1, 1, 35, 23, 1) op_2814 (v447[11:0], v1136[11:0], v2814[34:0]); // 3.0
    wire [23:0] v2815; shift_adder #(12, 21, 1, 1, 24, -11, 0) op_2815 (v1190[11:0], v1191[20:0], v2815[23:0]); // 3.0
    wire [34:0] v2816; shift_adder #(34, 22, 1, 1, 35, 12, 0) op_2816 (v1110[33:0], v1192[21:0], v2816[34:0]); // 3.0
    wire [13:0] v2817; shift_adder #(11, 14, 1, 1, 14, 0, 1) op_2817 (v232[10:0], v1002[13:0], v2817[13:0]); // 3.0
    wire [13:0] v2818; shift_adder #(13, 12, 1, 1, 14, 1, 0) op_2818 (v833[12:0], v239[11:0], v2818[13:0]); // 3.0
    wire [31:0] v2819; shift_adder #(32, 25, 1, 1, 32, 4, 0) op_2819 (v1193[31:0], v1194[24:0], v2819[31:0]); // 3.0
    wire [17:0] v2820; shift_adder #(11, 12, 1, 1, 18, 6, 0) op_2820 (v148[10:0], v971[11:0], v2820[17:0]); // 3.0
    wire [27:0] v2821; shift_adder #(13, 14, 1, 1, 28, -15, 0) op_2821 (v793[12:0], v1104[13:0], v2821[27:0]); // 3.0
    wire [21:0] v2822; shift_adder #(13, 19, 1, 1, 22, 3, 0) op_2822 (v449[12:0], v1195[18:0], v2822[21:0]); // 3.0
    wire [26:0] v2823; shift_adder #(8, 12, 1, 1, 27, 15, 1) op_2823 (v103[7:0], v1196[11:0], v2823[26:0]); // 3.0
    wire [28:0] v2824; shift_adder #(11, 21, 1, 1, 29, -18, 1) op_2824 (v418[10:0], v1197[20:0], v2824[28:0]); // 3.0
    wire [30:0] v2825; shift_adder #(12, 19, 1, 1, 31, -19, 1) op_2825 (v409[11:0], v1198[18:0], v2825[30:0]); // 3.0
    wire [22:0] v2826; shift_adder #(23, 16, 1, 1, 23, 5, 0) op_2826 (v1200[22:0], v1201[15:0], v2826[22:0]); // 3.0
    wire [24:0] v2827; shift_adder #(11, 13, 1, 1, 25, -14, 1) op_2827 (v157[10:0], v1202[12:0], v2827[24:0]); // 3.0
    wire [22:0] v2828; shift_adder #(12, 21, 1, 1, 23, -10, 0) op_2828 (v1203[11:0], v1128[20:0], v2828[22:0]); // 3.0
    wire [13:0] v2829; shift_adder #(11, 12, 1, 1, 14, 2, 0) op_2829 (v244[10:0], v981[11:0], v2829[13:0]); // 3.0
    wire [19:0] v2830; shift_adder #(16, 13, 1, 1, 20, 7, 0) op_2830 (v426[15:0], v845[12:0], v2830[19:0]); // 3.0
    wire [15:0] v2831; shift_adder #(14, 15, 1, 1, 16, 1, 0) op_2831 (v1204[13:0], v1205[14:0], v2831[15:0]); // 3.0
    wire [21:0] v2832; shift_adder #(12, 21, 1, 1, 22, -10, 1) op_2832 (v453[11:0], v1206[20:0], v2832[21:0]); // 3.0
    wire [29:0] v2833; shift_adder #(11, 25, 1, 1, 30, -19, 0) op_2833 (v455[10:0], v791[24:0], v2833[29:0]); // 3.0
    wire [19:0] v2834; shift_adder #(18, 18, 1, 1, 20, -1, 0) op_2834 (v1207[17:0], v1208[17:0], v2834[19:0]); // 3.0
    wire [17:0] v2835; shift_adder #(17, 17, 1, 1, 18, 1, 0) op_2835 (v852[16:0], v783[16:0], v2835[17:0]); // 3.0
    wire [12:0] v2836; shift_adder #(11, 13, 1, 1, 13, 0, 1) op_2836 (v145[10:0], v1209[12:0], v2836[12:0]); // 3.0
    wire [19:0] v2837; shift_adder #(19, 12, 1, 1, 20, 7, 0) op_2837 (v1210[18:0], v1211[11:0], v2837[19:0]); // 3.0
    wire [21:0] v2838; shift_adder #(21, 16, 1, 1, 22, 5, 0) op_2838 (v1212[20:0], v1213[15:0], v2838[21:0]); // 3.0
    wire [14:0] v2839; shift_adder #(11, 12, 1, 1, 15, 3, 0) op_2839 (v139[10:0], v1214[11:0], v2839[14:0]); // 3.0
    wire [25:0] v2840; shift_adder #(23, 21, 1, 1, 26, 5, 0) op_2840 (v1215[22:0], v1216[20:0], v2840[25:0]); // 3.0
    wire [20:0] v2841; shift_adder #(19, 19, 1, 1, 21, 2, 0) op_2841 (v1217[18:0], v1218[18:0], v2841[20:0]); // 3.0
    wire [28:0] v2842; shift_adder #(29, 17, 1, 1, 29, 11, 0) op_2842 (v1219[28:0], v1220[16:0], v2842[28:0]); // 3.0
    wire [21:0] v2843; shift_adder #(11, 17, 1, 1, 22, 5, 0) op_2843 (v1161[10:0], v1221[16:0], v2843[21:0]); // 3.0
    wire [29:0] v2844; shift_adder #(14, 30, 1, 1, 30, -15, 0) op_2844 (v1222[13:0], v1223[29:0], v2844[29:0]); // 3.0
    wire [20:0] v2845; shift_adder #(20, 15, 1, 1, 21, 5, 0) op_2845 (v1224[19:0], v1225[14:0], v2845[20:0]); // 3.0
    wire [20:0] v2846; shift_adder #(11, 19, 1, 1, 21, -10, 0) op_2846 (v455[10:0], v1226[18:0], v2846[20:0]); // 3.0
    wire [18:0] v2847; shift_adder #(11, 15, 1, 1, 19, 4, 1) op_2847 (v173[10:0], v1019[14:0], v2847[18:0]); // 3.0
    wire [13:0] v2848; shift_adder #(11, 13, 1, 1, 14, 1, 0) op_2848 (v297[10:0], v1079[12:0], v2848[13:0]); // 3.0
    wire [13:0] v2849; shift_adder #(12, 13, 1, 1, 14, 1, 0) op_2849 (v1004[11:0], v1227[12:0], v2849[13:0]); // 3.0
    wire [14:0] v2850; shift_adder #(14, 14, 1, 1, 15, 1, 0) op_2850 (v1228[13:0], v1229[13:0], v2850[14:0]); // 3.0
    wire [17:0] v2851; shift_adder #(10, 12, 1, 1, 18, -8, 0) op_2851 (v461[9:0], v1077[11:0], v2851[17:0]); // 3.0
    wire [21:0] v2852; shift_adder #(13, 17, 1, 1, 22, -9, 1) op_2852 (v1230[12:0], v1231[16:0], v2852[21:0]); // 3.0
    wire [29:0] v2853; shift_adder #(30, 14, 1, 1, 30, 15, 0) op_2853 (v1232[29:0], v1233[13:0], v2853[29:0]); // 3.0
    wire [24:0] v2854; shift_adder #(12, 23, 1, 1, 25, -13, 0) op_2854 (v1234[11:0], v1215[22:0], v2854[24:0]); // 3.0
    wire [20:0] v2855; shift_adder #(18, 17, 1, 1, 21, 4, 0) op_2855 (v1235[17:0], v1236[16:0], v2855[20:0]); // 3.0
    wire [23:0] v2856; shift_adder #(11, 19, 1, 1, 24, -13, 1) op_2856 (v241[10:0], v1237[18:0], v2856[23:0]); // 3.0
    wire [24:0] v2857; shift_adder #(13, 16, 1, 1, 25, -12, 0) op_2857 (v793[12:0], v1238[15:0], v2857[24:0]); // 3.0
    wire [30:0] v2858; shift_adder #(30, 11, 1, 1, 31, 19, 0) op_2858 (v1239[29:0], v1240[10:0], v2858[30:0]); // 3.0
    wire [15:0] v2859; shift_adder #(14, 12, 1, 1, 16, 3, 0) op_2859 (v1002[13:0], v1241[11:0], v2859[15:0]); // 3.0
    wire [12:0] v2860; shift_adder #(12, 13, 1, 1, 13, 0, 0) op_2860 (v288[11:0], v790[12:0], v2860[12:0]); // 3.0
    wire [28:0] v2861; shift_adder #(12, 28, 1, 1, 29, -17, 0) op_2861 (v1242[11:0], v1243[27:0], v2861[28:0]); // 3.0
    wire [21:0] v2862; shift_adder #(13, 10, 1, 1, 22, 12, 0) op_2862 (v1180[12:0], v470[9:0], v2862[21:0]); // 3.0
    wire [15:0] v2863; shift_adder #(8, 12, 1, 1, 16, 4, 1) op_2863 (v109[7:0], v1244[11:0], v2863[15:0]); // 3.0
    wire [28:0] v2864; shift_adder #(12, 28, 1, 1, 29, -16, 0) op_2864 (v990[11:0], v1245[27:0], v2864[28:0]); // 3.0
    wire [14:0] v2865; shift_adder #(13, 14, 1, 1, 15, 1, 0) op_2865 (v900[12:0], v472[13:0], v2865[14:0]); // 3.0
    wire [18:0] v2866; shift_adder #(19, 13, 1, 1, 19, 3, 1) op_2866 (v376[18:0], v995[12:0], v2866[18:0]); // 3.0
    wire [31:0] v2867; shift_adder #(8, 12, 1, 1, 32, -23, 1) op_2867 (v117[7:0], v896[11:0], v2867[31:0]); // 3.0
    wire [27:0] v2868; shift_adder #(27, 13, 1, 1, 28, 15, 0) op_2868 (v1246[26:0], v1247[12:0], v2868[27:0]); // 3.0
    wire [12:0] v2869; shift_adder #(8, 13, 1, 1, 13, -1, 0) op_2869 (v85[7:0], v1189[12:0], v2869[12:0]); // 3.0
    wire [16:0] v2870; shift_adder #(15, 16, 1, 1, 17, 0, 0) op_2870 (v1248[14:0], v1249[15:0], v2870[16:0]); // 3.0
    wire [13:0] v2871; shift_adder #(12, 14, 1, 1, 14, 0, 1) op_2871 (v292[11:0], v1250[13:0], v2871[13:0]); // 3.0
    wire [17:0] v2872; shift_adder #(14, 15, 1, 1, 18, -4, 0) op_2872 (v1251[13:0], v1252[14:0], v2872[17:0]); // 3.0
    wire [19:0] v2873; shift_adder #(9, 19, 1, 1, 20, -10, 1) op_2873 (v220[8:0], v944[18:0], v2873[19:0]); // 3.0
    wire [33:0] v2874; shift_adder #(13, 15, 1, 1, 34, -21, 1) op_2874 (v1041[12:0], v893[14:0], v2874[33:0]); // 3.0
    wire [16:0] v2875; shift_adder #(12, 15, 1, 1, 17, -5, 0) op_2875 (v1253[11:0], v1254[14:0], v2875[16:0]); // 3.0
    wire [12:0] v2876; shift_adder #(12, 12, 1, 1, 13, 0, 0) op_2876 (v365[11:0], v1255[11:0], v2876[12:0]); // 3.0
    wire [15:0] v2877; shift_adder #(14, 12, 1, 1, 16, 4, 0) op_2877 (v1256[13:0], v1257[11:0], v2877[15:0]); // 3.0
    wire [16:0] v2878; shift_adder #(12, 16, 1, 1, 17, -4, 0) op_2878 (v1258[11:0], v946[15:0], v2878[16:0]); // 3.0
    wire [12:0] v2879; shift_adder #(11, 12, 1, 1, 13, 1, 0) op_2879 (v455[10:0], v1259[11:0], v2879[12:0]); // 3.0
    wire [27:0] v2880; shift_adder #(27, 12, 1, 1, 28, 15, 0) op_2880 (v1260[26:0], v1261[11:0], v2880[27:0]); // 3.0
    wire [23:0] v2881; shift_adder #(12, 13, 1, 1, 24, -12, 1) op_2881 (v1262[11:0], v1263[12:0], v2881[23:0]); // 3.0
    wire [27:0] v2882; shift_adder #(9, 24, 1, 1, 28, 4, 1) op_2882 (v309[8:0], v1264[23:0], v2882[27:0]); // 3.0
    wire [28:0] v2883; shift_adder #(13, 15, 1, 1, 29, -16, 0) op_2883 (v813[12:0], v1265[14:0], v2883[28:0]); // 3.0
    wire [16:0] v2884; shift_adder #(17, 12, 1, 1, 17, 2, 0) op_2884 (v889[16:0], v1043[11:0], v2884[16:0]); // 3.0
    wire [20:0] v2885; shift_adder #(12, 21, 1, 1, 21, -7, 0) op_2885 (v423[11:0], v1266[20:0], v2885[20:0]); // 3.0
    wire [23:0] v2886; shift_adder #(21, 24, 1, 1, 24, -2, 0) op_2886 (v1267[20:0], v1268[23:0], v2886[23:0]); // 3.0
    wire [26:0] v2887; shift_adder #(25, 14, 1, 1, 27, 13, 0) op_2887 (v1269[24:0], v1270[13:0], v2887[26:0]); // 3.0
    wire [26:0] v2888; shift_adder #(27, 14, 1, 1, 27, 12, 0) op_2888 (v1271[26:0], v1112[13:0], v2888[26:0]); // 3.0
    wire [30:0] v2889; shift_adder #(8, 15, 1, 1, 31, 16, 1) op_2889 (v84[7:0], v1272[14:0], v2889[30:0]); // 3.0
    wire [28:0] v2890; shift_adder #(11, 27, 1, 1, 29, -18, 0) op_2890 (v1273[10:0], v1274[26:0], v2890[28:0]); // 3.0
    wire [16:0] v2891; shift_adder #(16, 12, 1, 1, 17, 4, 0) op_2891 (v1275[15:0], v1276[11:0], v2891[16:0]); // 3.0
    wire [12:0] v2892; shift_adder #(12, 12, 1, 1, 13, 0, 0) op_2892 (v1277[11:0], v1278[11:0], v2892[12:0]); // 3.0
    wire [14:0] v2893; shift_adder #(13, 13, 1, 1, 15, -2, 0) op_2893 (v859[12:0], v1279[12:0], v2893[14:0]); // 3.0
    wire [14:0] v2894; shift_adder #(8, 13, 1, 1, 15, 2, 1) op_2894 (v98[7:0], v1280[12:0], v2894[14:0]); // 3.0
    wire [15:0] v2895; shift_adder #(14, 15, 1, 1, 16, -1, 0) op_2895 (v1281[13:0], v1282[14:0], v2895[15:0]); // 3.0
    wire [12:0] v2896; shift_adder #(12, 11, 1, 1, 13, 0, 0) op_2896 (v1283[11:0], v1284[10:0], v2896[12:0]); // 3.0
    wire [20:0] v2897; shift_adder #(13, 15, 1, 1, 21, 6, 0) op_2897 (v1041[12:0], v1285[14:0], v2897[20:0]); // 3.0
    wire [24:0] v2898; shift_adder #(20, 24, 1, 1, 25, 1, 1) op_2898 (v1286[19:0], v1287[23:0], v2898[24:0]); // 3.0
    wire [23:0] v2899; shift_adder #(20, 14, 1, 1, 24, -4, 0) op_2899 (v484[19:0], v1288[13:0], v2899[23:0]); // 3.0
    wire [21:0] v2900; shift_adder #(8, 20, 1, 1, 22, 2, 0) op_2900 (v86[7:0], v1289[19:0], v2900[21:0]); // 3.0
    wire [13:0] v2901; shift_adder #(8, 14, 1, 1, 14, -3, 1) op_2901 (v102[7:0], v1290[13:0], v2901[13:0]); // 3.0
    wire [20:0] v2902; shift_adder #(17, 19, 1, 1, 21, -4, 0) op_2902 (v1291[16:0], v1292[18:0], v2902[20:0]); // 3.0
    wire [13:0] v2903; shift_adder #(11, 13, 1, 1, 14, -1, 0) op_2903 (v1293[10:0], v1294[12:0], v2903[13:0]); // 3.0
    wire [16:0] v2904; shift_adder #(13, 15, 1, 1, 17, -3, 0) op_2904 (v1295[12:0], v1296[14:0], v2904[16:0]); // 3.0
    wire [23:0] v2905; shift_adder #(23, 11, 1, 1, 24, 12, 0) op_2905 (v1297[22:0], v1298[10:0], v2905[23:0]); // 3.0
    wire [15:0] v2906; shift_adder #(14, 13, 1, 1, 16, 3, 0) op_2906 (v1299[13:0], v1163[12:0], v2906[15:0]); // 3.0
    wire [13:0] v2907; shift_adder #(11, 14, 1, 1, 14, 0, 0) op_2907 (v148[10:0], v1300[13:0], v2907[13:0]); // 3.0
    wire [13:0] v2908; shift_adder #(12, 14, 1, 1, 14, 0, 1) op_2908 (v265[11:0], v1301[13:0], v2908[13:0]); // 3.0
    wire [20:0] v2909; shift_adder #(8, 20, 1, 1, 21, 1, 1) op_2909 (v74[7:0], v1302[19:0], v2909[20:0]); // 3.0
    wire [15:0] v2910; shift_adder #(14, 15, 1, 1, 16, -1, 0) op_2910 (v1303[13:0], v1304[14:0], v2910[15:0]); // 3.0
    wire [17:0] v2911; shift_adder #(12, 11, 1, 1, 18, 7, 0) op_2911 (v1305[11:0], v1306[10:0], v2911[17:0]); // 3.0
    wire [14:0] v2912; shift_adder #(14, 12, 1, 1, 15, 3, 0) op_2912 (v1307[13:0], v1308[11:0], v2912[14:0]); // 3.0
    wire [22:0] v2913; shift_adder #(19, 22, 1, 1, 23, 1, 0) op_2913 (v805[18:0], v1179[21:0], v2913[22:0]); // 3.0
    wire [14:0] v2914; shift_adder #(12, 14, 1, 1, 15, -2, 1) op_2914 (v1309[11:0], v992[13:0], v2914[14:0]); // 3.0
    wire [22:0] v2915; shift_adder #(21, 14, 1, 1, 23, 9, 0) op_2915 (v1197[20:0], v1310[13:0], v2915[22:0]); // 3.0
    wire [15:0] v2916; shift_adder #(11, 16, 1, 1, 16, -4, 0) op_2916 (v139[10:0], v1311[15:0], v2916[15:0]); // 3.0
    wire [17:0] v2917; shift_adder #(17, 13, 1, 1, 18, 5, 0) op_2917 (v1312[16:0], v1029[12:0], v2917[17:0]); // 3.0
    wire [15:0] v2918; shift_adder #(9, 14, 1, 1, 16, -6, 1) op_2918 (v490[8:0], v1313[13:0], v2918[15:0]); // 3.0
    wire [17:0] v2919; shift_adder #(12, 17, 1, 1, 18, -5, 0) op_2919 (v1314[11:0], v1315[16:0], v2919[17:0]); // 3.0
    wire [16:0] v2920; shift_adder #(8, 13, 1, 1, 17, 4, 1) op_2920 (v89[7:0], v884[12:0], v2920[16:0]); // 3.0
    wire [17:0] v2921; shift_adder #(15, 18, 1, 1, 18, -2, 0) op_2921 (v840[14:0], v1316[17:0], v2921[17:0]); // 3.0
    wire [16:0] v2922; shift_adder #(14, 13, 1, 1, 17, 4, 0) op_2922 (v1317[13:0], v492[12:0], v2922[16:0]); // 3.0
    wire [32:0] v2923; shift_adder #(32, 13, 1, 1, 33, 19, 0) op_2923 (v1318[31:0], v892[12:0], v2923[32:0]); // 3.0
    wire [21:0] v2924; shift_adder #(11, 17, 1, 1, 22, -11, 1) op_2924 (v173[10:0], v783[16:0], v2924[21:0]); // 3.0
    wire [25:0] v2925; shift_adder #(13, 23, 1, 1, 26, 3, 1) op_2925 (v920[12:0], v1319[22:0], v2925[25:0]); // 3.0
    wire [27:0] v2926; shift_adder #(11, 19, 1, 1, 28, -17, 1) op_2926 (v375[10:0], v1320[18:0], v2926[27:0]); // 3.0
    wire [20:0] v2927; shift_adder #(19, 14, 1, 1, 21, 6, 0) op_2927 (v1321[18:0], v1162[13:0], v2927[20:0]); // 3.0
    wire [32:0] v2928; shift_adder #(11, 11, 1, 1, 33, 22, 1) op_2928 (v250[10:0], v885[10:0], v2928[32:0]); // 3.0
    wire [12:0] v2929; shift_adder #(11, 13, 1, 1, 13, -1, 1) op_2929 (v206[10:0], v1078[12:0], v2929[12:0]); // 3.0
    wire [32:0] v2930; shift_adder #(18, 33, 1, 1, 33, -1, 0) op_2930 (v493[17:0], v1322[32:0], v2930[32:0]); // 3.0
    wire [23:0] v2931; shift_adder #(19, 23, 1, 1, 24, -4, 0) op_2931 (v315[18:0], v1323[22:0], v2931[23:0]); // 3.0
    wire [16:0] v2932; shift_adder #(13, 15, 1, 1, 17, -4, 0) op_2932 (v1324[12:0], v781[14:0], v2932[16:0]); // 3.0
    wire [18:0] v2933; shift_adder #(18, 11, 1, 1, 19, 7, 0) op_2933 (v1325[17:0], v1137[10:0], v2933[18:0]); // 3.0
    wire [14:0] v2934; shift_adder #(13, 13, 1, 1, 15, 1, 0) op_2934 (v1326[12:0], v1327[12:0], v2934[14:0]); // 3.0
    wire [14:0] v2935; shift_adder #(13, 14, 1, 1, 15, -2, 0) op_2935 (v1328[12:0], v1329[13:0], v2935[14:0]); // 3.0
    wire [33:0] v2936; shift_adder #(15, 32, 1, 1, 34, -18, 0) op_2936 (v1330[14:0], v1331[31:0], v2936[33:0]); // 3.0
    wire [24:0] v2937; shift_adder #(11, 24, 1, 1, 25, -13, 0) op_2937 (v1161[10:0], v864[23:0], v2937[24:0]); // 3.0
    wire [15:0] v2938; shift_adder #(14, 12, 1, 1, 16, 3, 0) op_2938 (v1332[13:0], v1333[11:0], v2938[15:0]); // 3.0
    wire [12:0] v2939; shift_adder #(11, 11, 1, 1, 13, 2, 1) op_2939 (v772[10:0], v497[10:0], v2939[12:0]); // 3.0
    wire [21:0] v2940; shift_adder #(20, 22, 1, 1, 22, -1, 0) op_2940 (v1334[19:0], v1335[21:0], v2940[21:0]); // 3.0
    wire [24:0] v2941; shift_adder #(12, 13, 1, 1, 25, -13, 0) op_2941 (v452[11:0], v1336[12:0], v2941[24:0]); // 3.0
    wire [34:0] v2942; shift_adder #(34, 26, 1, 1, 35, 8, 0) op_2942 (v1337[33:0], v1338[25:0], v2942[34:0]); // 3.0
    wire [25:0] v2943; shift_adder #(25, 14, 1, 1, 26, 11, 0) op_2943 (v1095[24:0], v1339[13:0], v2943[25:0]); // 3.0
    wire [12:0] v2944; shift_adder #(8, 12, 1, 1, 13, -3, 1) op_2944 (v86[7:0], v1340[11:0], v2944[12:0]); // 3.0
    wire [24:0] v2945; shift_adder #(13, 17, 1, 1, 25, 8, 1) op_2945 (v149[12:0], v897[16:0], v2945[24:0]); // 3.0
    wire [28:0] v2946; shift_adder #(8, 21, 1, 1, 29, -20, 0) op_2946 (v112[7:0], v1062[20:0], v2946[28:0]); // 3.0
    wire [22:0] v2947; shift_adder #(17, 22, 1, 1, 23, -6, 0) op_2947 (v1341[16:0], v1342[21:0], v2947[22:0]); // 3.0
    wire [18:0] v2948; shift_adder #(11, 17, 1, 1, 19, -7, 0) op_2948 (v1298[10:0], v1343[16:0], v2948[18:0]); // 3.0
    wire [15:0] v2949; shift_adder #(11, 12, 1, 1, 16, -5, 0) op_2949 (v209[10:0], v971[11:0], v2949[15:0]); // 3.0
    wire [22:0] v2950; shift_adder #(19, 22, 1, 1, 23, -3, 0) op_2950 (v1344[18:0], v1345[21:0], v2950[22:0]); // 3.0
    wire [19:0] v2951; shift_adder #(11, 20, 1, 1, 20, -6, 0) op_2951 (v165[10:0], v925[19:0], v2951[19:0]); // 3.0
    wire [15:0] v2952; shift_adder #(11, 15, 1, 1, 16, -4, 0) op_2952 (v219[10:0], v1055[14:0], v2952[15:0]); // 3.0
    wire [13:0] v2953; shift_adder #(8, 13, 1, 1, 14, -5, 1) op_2953 (v116[7:0], v1346[12:0], v2953[13:0]); // 3.0
    wire [12:0] v2954; shift_adder #(12, 12, 1, 1, 13, 0, 0) op_2954 (v1347[11:0], v1348[11:0], v2954[12:0]); // 3.0
    wire [20:0] v2955; shift_adder #(13, 19, 1, 1, 21, -7, 0) op_2955 (v1349[12:0], v911[18:0], v2955[20:0]); // 3.0
    wire [12:0] v2956; shift_adder #(8, 13, 1, 1, 13, -2, 1) op_2956 (v96[7:0], v932[12:0], v2956[12:0]); // 3.0
    wire [16:0] v2957; shift_adder #(15, 15, 1, 1, 17, -2, 0) op_2957 (v1350[14:0], v1285[14:0], v2957[16:0]); // 3.0
    wire [14:0] v2958; shift_adder #(8, 15, 1, 1, 15, -5, 1) op_2958 (v126[7:0], v1351[14:0], v2958[14:0]); // 3.0
    wire [24:0] v2959; shift_adder #(15, 25, 1, 1, 25, -4, 1) op_2959 (v1352[14:0], v1194[24:0], v2959[24:0]); // 3.0
    wire [30:0] v2960; shift_adder #(22, 30, 1, 1, 31, -7, 0) op_2960 (v1353[21:0], v1354[29:0], v2960[30:0]); // 3.0
    wire [13:0] v2961; shift_adder #(14, 12, 1, 1, 14, 0, 1) op_2961 (v830[13:0], v1190[11:0], v2961[13:0]); // 3.0
    wire [24:0] v2962; shift_adder #(22, 13, 1, 1, 25, 12, 0) op_2962 (v1355[21:0], v1356[12:0], v2962[24:0]); // 3.0
    wire [14:0] v2963; shift_adder #(14, 11, 1, 1, 15, 3, 0) op_2963 (v1357[13:0], v1358[10:0], v2963[14:0]); // 3.0
    wire [29:0] v2964; shift_adder #(13, 29, 1, 1, 30, -16, 0) op_2964 (v1359[12:0], v1219[28:0], v2964[29:0]); // 3.0
    wire [12:0] v2965; shift_adder #(13, 9, 1, 1, 13, 0, 1) op_2965 (v1029[12:0], v368[8:0], v2965[12:0]); // 3.0
    wire [15:0] v2966; shift_adder #(16, 13, 1, 1, 16, 1, 0) op_2966 (v1360[15:0], v1361[12:0], v2966[15:0]); // 3.0
    wire [14:0] v2967; shift_adder #(11, 14, 1, 1, 15, -2, 0) op_2967 (v1362[10:0], v1332[13:0], v2967[14:0]); // 3.0
    wire [16:0] v2968; shift_adder #(11, 16, 1, 1, 17, -5, 0) op_2968 (v1363[10:0], v1364[15:0], v2968[16:0]); // 3.0
    wire [37:0] v2969; shift_adder #(22, 37, 1, 1, 38, -15, 0) op_2969 (v1365[21:0], v1366[36:0], v2969[37:0]); // 3.0
    wire [15:0] v2970; shift_adder #(8, 15, 1, 1, 16, -6, 1) op_2970 (v116[7:0], v1367[14:0], v2970[15:0]); // 3.0
    wire [30:0] v2971; shift_adder #(12, 30, 1, 1, 31, -17, 0) op_2971 (v1368[11:0], v1369[29:0], v2971[30:0]); // 3.0
    wire [17:0] v2972; shift_adder #(12, 16, 1, 1, 18, -5, 0) op_2972 (v1370[11:0], v1371[15:0], v2972[17:0]); // 3.0
    wire [11:0] v2973; shift_adder #(8, 12, 1, 1, 12, 0, 0) op_2973 (v70[7:0], v1372[11:0], v2973[11:0]); // 3.0
    wire [16:0] v2974; shift_adder #(12, 15, 1, 1, 17, -5, 0) op_2974 (v1373[11:0], v1374[14:0], v2974[16:0]); // 3.0
    wire [12:0] v2975; shift_adder #(8, 13, 1, 1, 13, -2, 1) op_2975 (v91[7:0], v1375[12:0], v2975[12:0]); // 3.0
    wire [14:0] v2976; shift_adder #(12, 14, 1, 1, 15, -2, 0) op_2976 (v1376[11:0], v1377[13:0], v2976[14:0]); // 3.0
    wire [15:0] v2977; shift_adder #(8, 14, 1, 1, 16, 2, 0) op_2977 (v101[7:0], v1378[13:0], v2977[15:0]); // 3.0
    wire [13:0] v2978; shift_adder #(13, 12, 1, 1, 14, 2, 0) op_2978 (v1030[12:0], v257[11:0], v2978[13:0]); // 3.0
    wire [14:0] v2979; shift_adder #(12, 14, 1, 1, 15, -1, 0) op_2979 (v1379[11:0], v1380[13:0], v2979[14:0]); // 3.0
    wire [15:0] v2980; shift_adder #(14, 16, 1, 1, 16, -1, 0) op_2980 (v1381[13:0], v1382[15:0], v2980[15:0]); // 3.0
    wire [19:0] v2981; shift_adder #(12, 20, 1, 1, 20, -7, 0) op_2981 (v1383[11:0], v1384[19:0], v2981[19:0]); // 3.0
    wire [14:0] v2982; shift_adder #(12, 13, 1, 1, 15, 2, 0) op_2982 (v355[11:0], v1385[12:0], v2982[14:0]); // 3.0
    wire [13:0] v2983; shift_adder #(13, 12, 1, 1, 14, 0, 0) op_2983 (v834[12:0], v500[11:0], v2983[13:0]); // 3.0
    wire [14:0] v2984; shift_adder #(13, 15, 1, 1, 15, -1, 0) op_2984 (v1079[12:0], v1012[14:0], v2984[14:0]); // 3.0
    wire [13:0] v2985; shift_adder #(11, 14, 1, 1, 14, -1, 1) op_2985 (v393[10:0], v1386[13:0], v2985[13:0]); // 3.0
    wire [16:0] v2986; shift_adder #(8, 17, 1, 1, 17, -2, 1) op_2986 (v122[7:0], v819[16:0], v2986[16:0]); // 3.0
    wire [14:0] v2987; shift_adder #(11, 12, 1, 1, 15, 3, 0) op_2987 (v162[10:0], v1047[11:0], v2987[14:0]); // 3.0
    wire [22:0] v2988; shift_adder #(15, 22, 1, 1, 23, -7, 0) op_2988 (v1387[14:0], v1388[21:0], v2988[22:0]); // 3.0
    wire [25:0] v2989; shift_adder #(16, 26, 1, 1, 26, -7, 0) op_2989 (v1389[15:0], v1390[25:0], v2989[25:0]); // 3.0
    wire [18:0] v2990; shift_adder #(18, 17, 1, 1, 19, 2, 0) op_2990 (v1391[17:0], v1392[16:0], v2990[18:0]); // 3.0
    wire [13:0] v2991; shift_adder #(13, 13, 1, 1, 14, 1, 0) op_2991 (v1393[12:0], v326[12:0], v2991[13:0]); // 3.0
    wire [15:0] v2992; shift_adder #(15, 12, 1, 1, 16, 4, 0) op_2992 (v1107[14:0], v1178[11:0], v2992[15:0]); // 3.0
    wire [21:0] v2993; shift_adder #(8, 14, 1, 1, 22, 8, 0) op_2993 (v123[7:0], v1394[13:0], v2993[21:0]); // 3.0
    wire [24:0] v2994; shift_adder #(11, 25, 1, 1, 25, -12, 0) op_2994 (v1395[10:0], v1396[24:0], v2994[24:0]); // 3.0
    wire [21:0] v2995; shift_adder #(13, 12, 1, 1, 22, -9, 1) op_2995 (v1397[12:0], v1398[11:0], v2995[21:0]); // 3.0
    wire [14:0] v2996; shift_adder #(12, 14, 1, 1, 15, -1, 0) op_2996 (v1399[11:0], v899[13:0], v2996[14:0]); // 3.0
    wire [21:0] v2997; shift_adder #(12, 20, 1, 1, 22, -10, 0) op_2997 (v174[11:0], v1400[19:0], v2997[21:0]); // 3.0
    wire [20:0] v2998; shift_adder #(8, 12, 1, 1, 21, -12, 1) op_2998 (v66[7:0], v801[11:0], v2998[20:0]); // 3.0
    wire [18:0] v2999; shift_adder #(12, 15, 1, 1, 19, 4, 1) op_2999 (v336[11:0], v1401[14:0], v2999[18:0]); // 3.0
    wire [15:0] v3000; shift_adder #(14, 16, 1, 1, 16, -1, 0) op_3000 (v1386[13:0], v1402[15:0], v3000[15:0]); // 3.0
    wire [21:0] v3001; shift_adder #(21, 13, 1, 1, 22, 9, 0) op_3001 (v1403[20:0], v932[12:0], v3001[21:0]); // 3.0
    wire [13:0] v3002; shift_adder #(11, 13, 1, 1, 14, -2, 1) op_3002 (v197[10:0], v1404[12:0], v3002[13:0]); // 3.0
    wire [30:0] v3003; shift_adder #(11, 25, 1, 1, 31, -20, 0) op_3003 (v386[10:0], v1405[24:0], v3003[30:0]); // 3.0
    wire [25:0] v3004; shift_adder #(13, 13, 1, 1, 26, 13, 0) op_3004 (v920[12:0], v1279[12:0], v3004[25:0]); // 3.0
    wire [25:0] v3005; shift_adder #(24, 17, 1, 1, 26, 9, 0) op_3005 (v1287[23:0], v1406[16:0], v3005[25:0]); // 3.0
    wire [16:0] v3006; shift_adder #(16, 16, 1, 1, 17, 1, 0) op_3006 (v1156[15:0], v1238[15:0], v3006[16:0]); // 3.0
    wire [21:0] v3007; shift_adder #(11, 13, 1, 1, 22, 9, 1) op_3007 (v294[10:0], v1407[12:0], v3007[21:0]); // 3.0
    wire [34:0] v3008; shift_adder #(12, 11, 1, 1, 35, -23, 1) op_3008 (v1408[11:0], v1409[10:0], v3008[34:0]); // 3.0
    wire [23:0] v3009; shift_adder #(18, 24, 1, 1, 24, -5, 0) op_3009 (v1235[17:0], v1149[23:0], v3009[23:0]); // 3.0
    wire [16:0] v3010; shift_adder #(17, 12, 1, 1, 17, 2, 0) op_3010 (v1410[16:0], v797[11:0], v3010[16:0]); // 3.0
    wire [19:0] v3011; shift_adder #(20, 12, 1, 1, 20, 7, 0) op_3011 (v1411[19:0], v1412[11:0], v3011[19:0]); // 3.0
    wire [16:0] v3012; shift_adder #(12, 16, 1, 1, 17, -5, 0) op_3012 (v1413[11:0], v1414[15:0], v3012[16:0]); // 3.0
    wire [13:0] v3013; shift_adder #(11, 13, 1, 1, 14, -2, 0) op_3013 (v1415[10:0], v1416[12:0], v3013[13:0]); // 3.0
    wire [23:0] v3014; shift_adder #(15, 24, 1, 1, 24, -1, 1) op_3014 (v1417[14:0], v1418[23:0], v3014[23:0]); // 3.0
    wire [12:0] v3015; shift_adder #(11, 12, 1, 1, 13, -1, 0) op_3015 (v1419[10:0], v835[11:0], v3015[12:0]); // 3.0
    wire [14:0] v3016; shift_adder #(13, 14, 1, 1, 15, -1, 0) op_3016 (v1397[12:0], v1420[13:0], v3016[14:0]); // 3.0
    wire [17:0] v3017; shift_adder #(17, 17, 1, 1, 18, -1, 0) op_3017 (v1315[16:0], v1221[16:0], v3017[17:0]); // 3.0
    wire [17:0] v3018; shift_adder #(11, 13, 1, 1, 18, 5, 0) op_3018 (v200[10:0], v1421[12:0], v3018[17:0]); // 3.0
    wire [15:0] v3019; shift_adder #(11, 13, 1, 1, 16, -5, 0) op_3019 (v136[10:0], v1422[12:0], v3019[15:0]); // 3.0
    wire [25:0] v3020; shift_adder #(11, 19, 1, 1, 26, -15, 0) op_3020 (v229[10:0], v1423[18:0], v3020[25:0]); // 3.0
    wire [19:0] v3021; shift_adder #(11, 13, 1, 1, 20, -9, 0) op_3021 (v269[10:0], v985[12:0], v3021[19:0]); // 3.0
    wire [33:0] v3022; shift_adder #(33, 16, 1, 1, 34, 17, 0) op_3022 (v1322[32:0], v1424[15:0], v3022[33:0]); // 3.0
    wire [19:0] v3023; shift_adder #(16, 11, 1, 1, 20, 9, 1) op_3023 (v1425[15:0], v1426[10:0], v3023[19:0]); // 3.0
    wire [12:0] v3024; shift_adder #(12, 11, 1, 1, 13, 1, 0) op_3024 (v820[11:0], v1427[10:0], v3024[12:0]); // 3.0
    wire [15:0] v3025; shift_adder #(15, 15, 1, 1, 16, 1, 1) op_3025 (v1429[14:0], v1430[14:0], v3025[15:0]); // 3.0
    wire [32:0] v3026; shift_adder #(13, 33, 1, 1, 33, -19, 0) op_3026 (v1431[12:0], v1432[32:0], v3026[32:0]); // 3.0
    wire [13:0] v3027; shift_adder #(13, 12, 1, 1, 14, 1, 0) op_3027 (v1433[12:0], v1000[11:0], v3027[13:0]); // 3.0
    wire [13:0] v3028; shift_adder #(10, 12, 1, 1, 14, -4, 0) op_3028 (v307[9:0], v1214[11:0], v3028[13:0]); // 3.0
    wire [37:0] v3029; shift_adder #(15, 37, 1, 1, 38, -22, 0) op_3029 (v1434[14:0], v1435[36:0], v3029[37:0]); // 3.0
    wire [13:0] v3030; shift_adder #(12, 12, 1, 1, 14, 1, 0) op_3030 (v1436[11:0], v1437[11:0], v3030[13:0]); // 3.0
    wire [14:0] v3031; shift_adder #(14, 13, 1, 1, 15, -1, 0) op_3031 (v1301[13:0], v1438[12:0], v3031[14:0]); // 3.0
    wire [14:0] v3032; shift_adder #(11, 15, 1, 1, 15, -1, 1) op_3032 (v250[10:0], v1439[14:0], v3032[14:0]); // 3.0
    wire [33:0] v3033; shift_adder #(13, 33, 1, 1, 34, -20, 0) op_3033 (v1440[12:0], v1441[32:0], v3033[33:0]); // 3.0
    wire [30:0] v3034; shift_adder #(30, 12, 1, 1, 31, 19, 0) op_3034 (v1442[29:0], v1443[11:0], v3034[30:0]); // 3.0
    wire [25:0] v3035; shift_adder #(25, 18, 1, 1, 26, 7, 0) op_3035 (v1444[24:0], v1445[17:0], v3035[25:0]); // 3.0
    wire [21:0] v3036; shift_adder #(11, 11, 1, 1, 22, -11, 1) op_3036 (v1161[10:0], v443[10:0], v3036[21:0]); // 3.0
    wire [21:0] v3037; shift_adder #(8, 13, 1, 1, 22, 9, 1) op_3037 (v99[7:0], v1446[12:0], v3037[21:0]); // 3.0
    wire [15:0] v3038; shift_adder #(8, 16, 1, 1, 16, -4, 1) op_3038 (v113[7:0], v1447[15:0], v3038[15:0]); // 3.0
    wire [26:0] v3039; shift_adder #(26, 26, 1, 1, 27, -1, 0) op_3039 (v1448[25:0], v1449[25:0], v3039[26:0]); // 3.0
    wire [23:0] v3040; shift_adder #(24, 12, 1, 1, 24, 10, 0) op_3040 (v1450[23:0], v1100[11:0], v3040[23:0]); // 3.0
    wire [26:0] v3041; shift_adder #(14, 26, 1, 1, 27, -12, 0) op_3041 (v1313[13:0], v1050[25:0], v3041[26:0]); // 3.0
    wire [17:0] v3042; shift_adder #(18, 16, 1, 1, 18, 1, 0) op_3042 (v1451[17:0], v1452[15:0], v3042[17:0]); // 3.0
    wire [25:0] v3043; shift_adder #(14, 18, 1, 1, 26, 8, 1) op_3043 (v481[13:0], v1453[17:0], v3043[25:0]); // 3.0
    wire [26:0] v3044; shift_adder #(26, 17, 1, 1, 27, 9, 0) op_3044 (v1454[25:0], v1455[16:0], v3044[26:0]); // 3.0
    wire [14:0] v3045; shift_adder #(9, 13, 1, 1, 15, -5, 0) op_3045 (v368[8:0], v900[12:0], v3045[14:0]); // 3.0
    wire [22:0] v3046; shift_adder #(13, 20, 1, 1, 23, -10, 0) op_3046 (v1456[12:0], v1457[19:0], v3046[22:0]); // 3.0
    wire [20:0] v3047; shift_adder #(13, 13, 1, 1, 21, -8, 0) op_3047 (v1458[12:0], v1459[12:0], v3047[20:0]); // 3.0
    wire [23:0] v3048; shift_adder #(11, 24, 1, 1, 24, -3, 0) op_3048 (v135[10:0], v1460[23:0], v3048[23:0]); // 3.0
    wire [13:0] v3049; shift_adder #(9, 13, 1, 1, 14, -3, 1) op_3049 (v531[8:0], v1461[12:0], v3049[13:0]); // 3.0
    wire [21:0] v3050; shift_adder #(12, 13, 1, 1, 22, -10, 0) op_3050 (v292[11:0], v813[12:0], v3050[21:0]); // 3.0
    wire [20:0] v3051; shift_adder #(8, 12, 1, 1, 21, -12, 1) op_3051 (v119[7:0], v1462[11:0], v3051[20:0]); // 3.0
    wire [23:0] v3052; shift_adder #(12, 21, 1, 1, 24, 3, 1) op_3052 (v862[11:0], v777[20:0], v3052[23:0]); // 3.0
    wire [12:0] v3053; shift_adder #(12, 13, 1, 1, 13, 0, 0) op_3053 (v1463[11:0], v1279[12:0], v3053[12:0]); // 3.0
    wire [16:0] v3054; shift_adder #(17, 11, 1, 1, 17, 5, 0) op_3054 (v1464[16:0], v1465[10:0], v3054[16:0]); // 3.0
    wire [19:0] v3055; shift_adder #(12, 20, 1, 1, 20, -6, 0) op_3055 (v1466[11:0], v809[19:0], v3055[19:0]); // 3.0
    wire [16:0] v3056; shift_adder #(17, 12, 1, 1, 17, 3, 0) op_3056 (v1467[16:0], v1468[11:0], v3056[16:0]); // 3.0
    wire [23:0] v3057; shift_adder #(23, 24, 1, 1, 24, 0, 0) op_3057 (v1469[22:0], v1470[23:0], v3057[23:0]); // 3.0
    wire [15:0] v3058; shift_adder #(13, 16, 1, 1, 16, -1, 0) op_3058 (v1471[12:0], v1472[15:0], v3058[15:0]); // 3.0
    wire [19:0] v3059; shift_adder #(13, 13, 1, 1, 20, -7, 1) op_3059 (v1029[12:0], v884[12:0], v3059[19:0]); // 3.0
    wire [23:0] v3060; shift_adder #(15, 12, 1, 1, 24, 12, 0) op_3060 (v1473[14:0], v532[11:0], v3060[23:0]); // 3.0
    wire [13:0] v3061; shift_adder #(8, 13, 1, 1, 14, -4, 0) op_3061 (v68[7:0], v891[12:0], v3061[13:0]); // 3.0
    wire [22:0] v3062; shift_adder #(16, 23, 1, 1, 23, -6, 0) op_3062 (v1089[15:0], v1474[22:0], v3062[22:0]); // 3.0
    wire [21:0] v3063; shift_adder #(22, 14, 1, 1, 22, 7, 0) op_3063 (v774[21:0], v1072[13:0], v3063[21:0]); // 3.0
    wire [26:0] v3064; shift_adder #(12, 27, 1, 1, 27, -14, 0) op_3064 (v1475[11:0], v1476[26:0], v3064[26:0]); // 3.0
    wire [16:0] v3065; shift_adder #(12, 17, 1, 1, 17, -4, 0) op_3065 (v973[11:0], v967[16:0], v3065[16:0]); // 3.0
    wire [19:0] v3066; shift_adder #(8, 15, 1, 1, 20, 5, 1) op_3066 (v113[7:0], v1477[14:0], v3066[19:0]); // 3.0
    wire [17:0] v3067; shift_adder #(17, 13, 1, 1, 18, 4, 0) op_3067 (v1478[16:0], v1479[12:0], v3067[17:0]); // 3.0
    wire [17:0] v3068; shift_adder #(13, 18, 1, 1, 18, -4, 0) op_3068 (v915[12:0], v535[17:0], v3068[17:0]); // 3.0
    wire [19:0] v3069; shift_adder #(14, 20, 1, 1, 20, -4, 0) op_3069 (v1480[13:0], v1481[19:0], v3069[19:0]); // 3.0
    wire [27:0] v3070; shift_adder #(10, 13, 1, 1, 28, 15, 0) op_3070 (v469[9:0], v1482[12:0], v3070[27:0]); // 3.0
    wire [31:0] v3071; shift_adder #(31, 30, 1, 1, 32, -1, 0) op_3071 (v1140[30:0], v1354[29:0], v3071[31:0]); // 3.0
    wire [21:0] v3072; shift_adder #(14, 12, 1, 1, 22, -8, 0) op_3072 (v1307[13:0], v1103[11:0], v3072[21:0]); // 3.0
    wire [25:0] v3073; shift_adder #(16, 26, 1, 1, 26, -7, 0) op_3073 (v1213[15:0], v1483[25:0], v3073[25:0]); // 3.0
    wire [17:0] v3074; shift_adder #(14, 12, 1, 1, 18, 6, 0) op_3074 (v1250[13:0], v1484[11:0], v3074[17:0]); // 3.0
    wire [26:0] v3075; shift_adder #(17, 26, 1, 1, 27, -9, 0) op_3075 (v1485[16:0], v1486[25:0], v3075[26:0]); // 3.0
    wire [31:0] v3076; shift_adder #(13, 24, 1, 1, 32, -19, 1) op_3076 (v492[12:0], v1487[23:0], v3076[31:0]); // 3.0
    wire [26:0] v3077; shift_adder #(8, 14, 1, 1, 27, -18, 1) op_3077 (v76[7:0], v975[13:0], v3077[26:0]); // 3.0
    wire [31:0] v3078; shift_adder #(31, 25, 1, 1, 32, 7, 0) op_3078 (v1488[30:0], v1092[24:0], v3078[31:0]); // 3.0
    wire [23:0] v3079; shift_adder #(13, 16, 1, 1, 24, -11, 0) op_3079 (v1397[12:0], v1238[15:0], v3079[23:0]); // 3.0
    wire [35:0] v3080; shift_adder #(36, 13, 1, 1, 36, 0, 1) op_3080 (v1489[35:0], v1490[12:0], v3080[35:0]); // 3.0
    wire [37:0] v3081; shift_adder #(13, 10, 1, 1, 38, 28, 1) op_3081 (v1189[12:0], v520[9:0], v3081[37:0]); // 3.0
    wire [12:0] v3082; shift_adder #(12, 11, 1, 1, 13, 1, 0) op_3082 (v1491[11:0], v1492[10:0], v3082[12:0]); // 3.0
    wire [12:0] v3083; shift_adder #(12, 9, 1, 1, 13, 1, 1) op_3083 (v1493[11:0], v467[8:0], v3083[12:0]); // 3.0
    wire [12:0] v3084; shift_adder #(11, 13, 1, 1, 13, -1, 0) op_3084 (v1494[10:0], v1495[12:0], v3084[12:0]); // 3.0
    wire [14:0] v3085; shift_adder #(14, 13, 1, 1, 15, 1, 0) op_3085 (v1496[13:0], v1497[12:0], v3085[14:0]); // 3.0
    wire [14:0] v3086; shift_adder #(14, 12, 1, 1, 15, 2, 0) op_3086 (v1126[13:0], v1498[11:0], v3086[14:0]); // 3.0
    wire [15:0] v3087; shift_adder #(15, 11, 1, 1, 16, 4, 0) op_3087 (v1499[14:0], v855[10:0], v3087[15:0]); // 3.0
    wire [13:0] v3088; shift_adder #(13, 12, 1, 1, 14, 1, 0) op_3088 (v1500[12:0], v1155[11:0], v3088[13:0]); // 3.0
    wire [18:0] v3089; shift_adder #(13, 18, 1, 1, 19, -5, 0) op_3089 (v1501[12:0], v1502[17:0], v3089[18:0]); // 3.0
    wire [28:0] v3090; shift_adder #(16, 28, 1, 1, 29, -12, 0) op_3090 (v1503[15:0], v1504[27:0], v3090[28:0]); // 3.0
    wire [15:0] v3091; shift_adder #(13, 13, 1, 1, 16, -3, 0) op_3091 (v1030[12:0], v834[12:0], v3091[15:0]); // 3.0
    wire [20:0] v3092; shift_adder #(20, 13, 1, 1, 21, 7, 0) op_3092 (v1457[19:0], v1086[12:0], v3092[20:0]); // 3.0
    wire [12:0] v3093; shift_adder #(10, 13, 1, 1, 13, 0, 0) op_3093 (v282[9:0], v1375[12:0], v3093[12:0]); // 3.0
    wire [18:0] v3094; shift_adder #(19, 12, 1, 1, 19, 2, 0) op_3094 (v1505[18:0], v1506[11:0], v3094[18:0]); // 3.0
    wire [14:0] v3095; shift_adder #(14, 13, 1, 1, 15, 0, 0) op_3095 (v1507[13:0], v1508[12:0], v3095[14:0]); // 3.0
    wire [13:0] v3096; shift_adder #(8, 14, 1, 1, 14, -2, 0) op_3096 (v93[7:0], v1509[13:0], v3096[13:0]); // 3.0
    wire [17:0] v3097; shift_adder #(8, 18, 1, 1, 18, -3, 1) op_3097 (v90[7:0], v1510[17:0], v3097[17:0]); // 3.0
    wire [18:0] v3098; shift_adder #(12, 17, 1, 1, 19, -6, 0) op_3098 (v1511[11:0], v1455[16:0], v3098[18:0]); // 3.0
    wire [25:0] v3099; shift_adder #(11, 13, 1, 1, 26, 13, 0) op_3099 (v175[10:0], v1030[12:0], v3099[25:0]); // 3.0
    wire [11:0] v3100; shift_adder #(8, 12, 1, 1, 12, 0, 0) op_3100 (v95[7:0], v1512[11:0], v3100[11:0]); // 3.0
    wire [14:0] v3101; shift_adder #(13, 14, 1, 1, 15, -1, 0) op_3101 (v826[12:0], v786[13:0], v3101[14:0]); // 3.0
    wire [14:0] v3102; shift_adder #(14, 12, 1, 1, 15, 1, 0) op_3102 (v1513[13:0], v1514[11:0], v3102[14:0]); // 3.0
    wire [19:0] v3103; shift_adder #(11, 17, 1, 1, 20, -8, 0) op_3103 (v1122[10:0], v1016[16:0], v3103[19:0]); // 3.0
    wire [23:0] v3104; shift_adder #(12, 24, 1, 1, 24, -1, 0) op_3104 (v550[11:0], v1515[23:0], v3104[23:0]); // 3.0
    wire [14:0] v3105; shift_adder #(11, 14, 1, 1, 15, -3, 0) op_3105 (v393[10:0], v1516[13:0], v3105[14:0]); // 3.0
    wire [13:0] v3106; shift_adder #(14, 12, 1, 1, 14, 1, 1) op_3106 (v1307[13:0], v354[11:0], v3106[13:0]); // 3.0
    wire [12:0] v3107; shift_adder #(9, 11, 1, 1, 13, -3, 0) op_3107 (v433[8:0], v1517[10:0], v3107[12:0]); // 3.0
    wire [17:0] v3108; shift_adder #(13, 17, 1, 1, 18, -4, 0) op_3108 (v1518[12:0], v1519[16:0], v3108[17:0]); // 3.0
    wire [20:0] v3109; shift_adder #(11, 13, 1, 1, 21, -10, 1) op_3109 (v197[10:0], v1421[12:0], v3109[20:0]); // 3.0
    wire [21:0] v3110; shift_adder #(21, 12, 1, 1, 22, 10, 0) op_3110 (v1520[20:0], v1521[11:0], v3110[21:0]); // 3.0
    wire [15:0] v3111; shift_adder #(14, 13, 1, 1, 16, 2, 0) op_3111 (v1522[13:0], v1349[12:0], v3111[15:0]); // 3.0
    wire [15:0] v3112; shift_adder #(11, 16, 1, 1, 16, -3, 0) op_3112 (v1523[10:0], v1311[15:0], v3112[15:0]); // 3.0
    wire [20:0] v3113; shift_adder #(19, 14, 1, 1, 21, 7, 0) op_3113 (v1113[18:0], v1303[13:0], v3113[20:0]); // 3.0
    wire [14:0] v3114; shift_adder #(14, 14, 1, 1, 15, 0, 0) op_3114 (v1039[13:0], v1303[13:0], v3114[14:0]); // 3.0
    wire [23:0] v3115; shift_adder #(11, 13, 1, 1, 24, 11, 0) op_3115 (v157[10:0], v1524[12:0], v3115[23:0]); // 3.0
    wire [28:0] v3116; shift_adder #(16, 17, 1, 1, 29, 12, 1) op_3116 (v1525[15:0], v1526[16:0], v3116[28:0]); // 3.0
    wire [18:0] v3117; shift_adder #(13, 19, 1, 1, 19, -5, 1) op_3117 (v1336[12:0], v1527[18:0], v3117[18:0]); // 3.0
    wire [27:0] v3118; shift_adder #(28, 17, 1, 1, 28, 10, 0) op_3118 (v1528[27:0], v773[16:0], v3118[27:0]); // 3.0
    wire [12:0] v3119; shift_adder #(9, 12, 1, 1, 13, -3, 0) op_3119 (v531[8:0], v1529[11:0], v3119[12:0]); // 3.0
    wire [25:0] v3120; shift_adder #(12, 19, 1, 1, 26, 7, 0) op_3120 (v553[11:0], v1530[18:0], v3120[25:0]); // 3.0
    wire [23:0] v3121; shift_adder #(8, 16, 1, 1, 24, -15, 1) op_3121 (v94[7:0], v1531[15:0], v3121[23:0]); // 3.0
    wire [14:0] v3122; shift_adder #(14, 13, 1, 1, 15, 0, 0) op_3122 (v1532[13:0], v1533[12:0], v3122[14:0]); // 3.0
    wire [22:0] v3123; shift_adder #(12, 12, 1, 1, 23, -11, 1) op_3123 (v453[11:0], v1534[11:0], v3123[22:0]); // 3.0
    wire [15:0] v3124; shift_adder #(15, 15, 1, 1, 16, -1, 1) op_3124 (v1535[14:0], v1536[14:0], v3124[15:0]); // 3.0
    wire [16:0] v3125; shift_adder #(12, 14, 1, 1, 17, 3, 1) op_3125 (v1537[11:0], v1538[13:0], v3125[16:0]); // 3.0
    wire [21:0] v3126; shift_adder #(13, 21, 1, 1, 22, -9, 0) op_3126 (v1187[12:0], v1539[20:0], v3126[21:0]); // 3.0
    wire [27:0] v3127; shift_adder #(11, 17, 1, 1, 28, 11, 1) op_3127 (v145[10:0], v1540[16:0], v3127[27:0]); // 3.0
    wire [17:0] v3128; shift_adder #(15, 16, 1, 1, 18, -3, 0) op_3128 (v969[14:0], v1106[15:0], v3128[17:0]); // 3.0
    wire [17:0] v3129; shift_adder #(16, 16, 1, 1, 18, -2, 0) op_3129 (v426[15:0], v1541[15:0], v3129[17:0]); // 3.0
    wire [17:0] v3130; shift_adder #(16, 17, 1, 1, 18, 1, 0) op_3130 (v1156[15:0], v1542[16:0], v3130[17:0]); // 3.0
    wire [17:0] v3131; shift_adder #(13, 14, 1, 1, 18, 4, 0) op_3131 (v883[12:0], v1538[13:0], v3131[17:0]); // 3.0
    wire [20:0] v3132; shift_adder #(18, 11, 1, 1, 21, 10, 0) op_3132 (v1096[17:0], v1543[10:0], v3132[20:0]); // 3.0
    wire [24:0] v3133; shift_adder #(8, 11, 1, 1, 25, 14, 0) op_3133 (v73[7:0], v846[10:0], v3133[24:0]); // 3.0
    wire [24:0] v3134; shift_adder #(14, 25, 1, 1, 25, -9, 0) op_3134 (v226[13:0], v1544[24:0], v3134[24:0]); // 3.0
    wire [13:0] v3135; shift_adder #(8, 11, 1, 1, 14, -5, 0) op_3135 (v74[7:0], v821[10:0], v3135[13:0]); // 3.0
    wire [13:0] v3136; shift_adder #(12, 14, 1, 1, 14, 0, 0) op_3136 (v457[11:0], v1545[13:0], v3136[13:0]); // 3.0
    wire [19:0] v3137; shift_adder #(17, 19, 1, 1, 20, -2, 0) op_3137 (v1546[16:0], v1547[18:0], v3137[19:0]); // 3.0
    wire [22:0] v3138; shift_adder #(11, 12, 1, 1, 23, -12, 0) op_3138 (v190[10:0], v1534[11:0], v3138[22:0]); // 3.0
    wire [23:0] v3139; shift_adder #(24, 17, 1, 1, 24, 6, 0) op_3139 (v1548[23:0], v881[16:0], v3139[23:0]); // 3.0
    wire [13:0] v3140; shift_adder #(14, 12, 1, 1, 14, 0, 0) op_3140 (v1549[13:0], v1550[11:0], v3140[13:0]); // 3.0
    wire [18:0] v3141; shift_adder #(13, 17, 1, 1, 19, -5, 0) op_3141 (v1551[12:0], v982[16:0], v3141[18:0]); // 3.0
    wire [16:0] v3142; shift_adder #(14, 16, 1, 1, 17, -3, 0) op_3142 (v799[13:0], v1552[15:0], v3142[16:0]); // 3.0
    wire [18:0] v3143; shift_adder #(19, 14, 1, 1, 19, 4, 0) op_3143 (v1553[18:0], v1554[13:0], v3143[18:0]); // 3.0
    wire [20:0] v3144; shift_adder #(21, 12, 1, 1, 21, 7, 0) op_3144 (v1040[20:0], v808[11:0], v3144[20:0]); // 3.0
    wire [18:0] v3145; shift_adder #(11, 12, 1, 1, 19, -8, 1) op_3145 (v238[10:0], v1555[11:0], v3145[18:0]); // 3.0
    wire [14:0] v3146; shift_adder #(12, 12, 1, 1, 15, -3, 0) op_3146 (v1379[11:0], v1556[11:0], v3146[14:0]); // 3.0
    wire [20:0] v3147; shift_adder #(11, 16, 1, 1, 21, -10, 1) op_3147 (v175[10:0], v1557[15:0], v3147[20:0]); // 3.0
    wire [13:0] v3148; shift_adder #(12, 13, 1, 1, 14, -2, 0) op_3148 (v1558[11:0], v1559[12:0], v3148[13:0]); // 3.0
    wire [13:0] v3149; shift_adder #(9, 13, 1, 1, 14, -3, 1) op_3149 (v368[8:0], v1560[12:0], v3149[13:0]); // 3.0
    wire [24:0] v3150; shift_adder #(18, 24, 1, 1, 25, -6, 0) op_3150 (v1561[17:0], v1460[23:0], v3150[24:0]); // 3.0
    wire [12:0] v3151; shift_adder #(8, 13, 1, 1, 13, -3, 0) op_3151 (v86[7:0], v1397[12:0], v3151[12:0]); // 3.0
    wire [16:0] v3152; shift_adder #(11, 12, 1, 1, 17, -6, 0) op_3152 (v216[10:0], v794[11:0], v3152[16:0]); // 3.0
    wire [21:0] v3153; shift_adder #(22, 12, 1, 1, 22, 8, 0) op_3153 (v1562[21:0], v1277[11:0], v3153[21:0]); // 3.0
    wire [18:0] v3154; shift_adder #(15, 18, 1, 1, 19, -4, 0) op_3154 (v914[14:0], v1563[17:0], v3154[18:0]); // 3.0
    wire [17:0] v3155; shift_adder #(18, 16, 1, 1, 18, 0, 0) op_3155 (v1099[17:0], v1564[15:0], v3155[17:0]); // 3.0
    wire [19:0] v3156; shift_adder #(13, 19, 1, 1, 20, -7, 0) op_3156 (v880[12:0], v1226[18:0], v3156[19:0]); // 3.0
    wire [12:0] v3157; shift_adder #(8, 13, 1, 1, 13, -1, 1) op_3157 (v65[7:0], v859[12:0], v3157[12:0]); // 3.0
    wire [19:0] v3158; shift_adder #(12, 19, 1, 1, 20, -7, 0) op_3158 (v434[11:0], v1565[18:0], v3158[19:0]); // 3.0
    wire [14:0] v3159; shift_adder #(12, 11, 1, 1, 15, -3, 0) op_3159 (v1566[11:0], v1298[10:0], v3159[14:0]); // 3.0
    wire [21:0] v3160; shift_adder #(20, 19, 1, 1, 22, 3, 0) op_3160 (v1567[19:0], v1568[18:0], v3160[21:0]); // 3.0
    wire [22:0] v3161; shift_adder #(8, 13, 1, 1, 23, 10, 1) op_3161 (v106[7:0], v1569[12:0], v3161[22:0]); // 3.0
    wire [19:0] v3162; shift_adder #(17, 15, 1, 1, 20, 4, 0) op_3162 (v1343[16:0], v1330[14:0], v3162[19:0]); // 3.0
    wire [19:0] v3163; shift_adder #(8, 12, 1, 1, 20, 8, 0) op_3163 (v95[7:0], v1570[11:0], v3163[19:0]); // 3.0
    wire [17:0] v3164; shift_adder #(14, 12, 1, 1, 18, -4, 0) op_3164 (v290[13:0], v1571[11:0], v3164[17:0]); // 3.0
    wire [15:0] v3165; shift_adder #(8, 15, 1, 1, 16, -6, 1) op_3165 (v108[7:0], v1572[14:0], v3165[15:0]); // 3.0
    wire [20:0] v3166; shift_adder #(8, 12, 1, 1, 21, 9, 0) op_3166 (v86[7:0], v1573[11:0], v3166[20:0]); // 3.0
    wire [19:0] v3167; shift_adder #(17, 14, 1, 1, 20, 6, 0) op_3167 (v1574[16:0], v1575[13:0], v3167[19:0]); // 3.0
    wire [22:0] v3168; shift_adder #(8, 13, 1, 1, 23, -14, 1) op_3168 (v109[7:0], v1079[12:0], v3168[22:0]); // 3.0
    wire [15:0] v3169; shift_adder #(11, 15, 1, 1, 16, -4, 0) op_3169 (v195[10:0], v1576[14:0], v3169[15:0]); // 3.0
    wire [15:0] v3170; shift_adder #(13, 15, 1, 1, 16, -2, 0) op_3170 (v828[12:0], v1577[14:0], v3170[15:0]); // 3.0
    wire [23:0] v3171; shift_adder #(24, 16, 1, 1, 24, 6, 0) op_3171 (v1578[23:0], v1531[15:0], v3171[23:0]); // 3.0
    wire [26:0] v3172; shift_adder #(27, 23, 1, 1, 27, 3, 0) op_3172 (v1579[26:0], v1200[22:0], v3172[26:0]); // 3.0
    wire [19:0] v3173; shift_adder #(13, 20, 1, 1, 20, -5, 0) op_3173 (v932[12:0], v1580[19:0], v3173[19:0]); // 3.0
    wire [11:0] v3174; shift_adder #(10, 11, 1, 1, 12, -1, 1) op_3174 (v263[9:0], v1581[10:0], v3174[11:0]); // 3.0
    wire [25:0] v3175; shift_adder #(12, 26, 1, 1, 26, -12, 0) op_3175 (v801[11:0], v802[25:0], v3175[25:0]); // 3.0
    wire [22:0] v3176; shift_adder #(11, 13, 1, 1, 23, -12, 1) op_3176 (v418[10:0], v1034[12:0], v3176[22:0]); // 3.0
    wire [15:0] v3177; shift_adder #(13, 16, 1, 1, 16, -1, 0) op_3177 (v1582[12:0], v1311[15:0], v3177[15:0]); // 3.0
    wire [19:0] v3178; shift_adder #(11, 16, 1, 1, 20, -9, 1) op_3178 (v358[10:0], v1213[15:0], v3178[19:0]); // 3.0
    wire [16:0] v3179; shift_adder #(16, 16, 1, 1, 17, 0, 0) op_3179 (v1238[15:0], v350[15:0], v3179[16:0]); // 3.0
    wire [16:0] v3180; shift_adder #(15, 12, 1, 1, 17, 4, 0) op_3180 (v1583[14:0], v1584[11:0], v3180[16:0]); // 3.0
    wire [16:0] v3181; shift_adder #(12, 14, 1, 1, 17, 3, 0) op_3181 (v1585[11:0], v871[13:0], v3181[16:0]); // 3.0
    wire [21:0] v3182; shift_adder #(21, 16, 1, 1, 22, 5, 0) op_3182 (v1586[20:0], v1587[15:0], v3182[21:0]); // 3.0
    wire [22:0] v3183; shift_adder #(17, 23, 1, 1, 23, 0, 0) op_3183 (v1151[16:0], v1469[22:0], v3183[22:0]); // 3.0
    wire [26:0] v3184; shift_adder #(15, 13, 1, 1, 27, -12, 0) op_3184 (v1015[14:0], v1588[12:0], v3184[26:0]); // 3.0
    wire [28:0] v3185; shift_adder #(12, 9, 1, 1, 29, 19, 0) op_3185 (v1589[11:0], v477[8:0], v3185[28:0]); // 3.0
    wire [14:0] v3186; shift_adder #(8, 15, 1, 1, 15, -5, 1) op_3186 (v76[7:0], v1590[14:0], v3186[14:0]); // 3.0
    wire [17:0] v3187; shift_adder #(13, 18, 1, 1, 18, -3, 0) op_3187 (v1591[12:0], v1592[17:0], v3187[17:0]); // 3.0
    wire [19:0] v3188; shift_adder #(19, 13, 1, 1, 20, 7, 0) op_3188 (v1593[18:0], v1594[12:0], v3188[19:0]); // 3.0
    wire [30:0] v3189; shift_adder #(12, 16, 1, 1, 31, -19, 0) op_3189 (v553[11:0], v1552[15:0], v3189[30:0]); // 3.0
    wire [22:0] v3190; shift_adder #(11, 23, 1, 1, 23, -10, 0) op_3190 (v962[10:0], v1595[22:0], v3190[22:0]); // 3.0
    wire [27:0] v3191; shift_adder #(21, 14, 1, 1, 28, -7, 1) op_3191 (v1596[20:0], v1513[13:0], v3191[27:0]); // 3.0
    wire [37:0] v3192; shift_adder #(34, 38, 1, 1, 38, -3, 0) op_3192 (v1597[33:0], v1598[37:0], v3192[37:0]); // 3.0
    wire [33:0] v3193; shift_adder #(13, 10, 1, 1, 34, 24, 1) op_3193 (v1599[12:0], v565[9:0], v3193[33:0]); // 3.0
    wire [13:0] v3194; shift_adder #(13, 12, 1, 1, 14, 0, 0) op_3194 (v817[12:0], v1600[11:0], v3194[13:0]); // 3.0
    wire [23:0] v3195; shift_adder #(12, 13, 1, 1, 24, 11, 1) op_3195 (v473[11:0], v837[12:0], v3195[23:0]); // 3.0
    wire [15:0] v3196; shift_adder #(12, 14, 1, 1, 16, -3, 0) op_3196 (v1602[11:0], v1299[13:0], v3196[15:0]); // 3.0
    wire [38:0] v3197; shift_adder #(20, 12, 1, 1, 39, -19, 1) op_3197 (v1603[19:0], v1604[11:0], v3197[38:0]); // 3.0
    wire [21:0] v3198; shift_adder #(20, 12, 1, 1, 22, 9, 0) op_3198 (v925[19:0], v1605[11:0], v3198[21:0]); // 3.0
    wire [17:0] v3199; shift_adder #(16, 13, 1, 1, 18, 4, 0) op_3199 (v1606[15:0], v920[12:0], v3199[17:0]); // 3.0
    wire [13:0] v3200; shift_adder #(14, 13, 1, 1, 14, 0, 0) op_3200 (v1607[13:0], v996[12:0], v3200[13:0]); // 3.0
    wire [14:0] v3201; shift_adder #(13, 13, 1, 1, 15, -2, 0) op_3201 (v880[12:0], v1608[12:0], v3201[14:0]); // 3.0
    wire [14:0] v3202; shift_adder #(15, 11, 1, 1, 15, 2, 0) op_3202 (v1609[14:0], v846[10:0], v3202[14:0]); // 3.0
    wire [17:0] v3203; shift_adder #(14, 15, 1, 1, 18, 3, 0) op_3203 (v1610[13:0], v1611[14:0], v3203[17:0]); // 3.0
    wire [13:0] v3204; shift_adder #(12, 12, 1, 1, 14, 1, 0) op_3204 (v1153[11:0], v1612[11:0], v3204[13:0]); // 3.0
    wire [15:0] v3205; shift_adder #(8, 11, 1, 1, 16, -7, 1) op_3205 (v104[7:0], v1613[10:0], v3205[15:0]); // 3.0
    wire [13:0] v3206; shift_adder #(12, 11, 1, 1, 14, 2, 0) op_3206 (v1614[11:0], v1615[10:0], v3206[13:0]); // 3.0
    wire [15:0] v3207; shift_adder #(11, 15, 1, 1, 16, 1, 0) op_3207 (v298[10:0], v839[14:0], v3207[15:0]); // 3.0
    wire [17:0] v3208; shift_adder #(13, 17, 1, 1, 18, -3, 0) op_3208 (v1616[12:0], v1617[16:0], v3208[17:0]); // 3.0
    wire [17:0] v3209; shift_adder #(17, 17, 1, 1, 18, 1, 0) op_3209 (v1618[16:0], v1619[16:0], v3209[17:0]); // 3.0
    wire [22:0] v3210; shift_adder #(16, 16, 1, 1, 23, 7, 1) op_3210 (v1620[15:0], v778[15:0], v3210[22:0]); // 3.0
    wire [25:0] v3211; shift_adder #(25, 13, 1, 1, 26, 12, 0) op_3211 (v1544[24:0], v1621[12:0], v3211[25:0]); // 3.0
    wire [23:0] v3212; shift_adder #(12, 24, 1, 1, 24, -2, 1) op_3212 (v1534[11:0], v1622[23:0], v3212[23:0]); // 3.0
    wire [17:0] v3213; shift_adder #(14, 17, 1, 1, 18, 1, 0) op_3213 (v1623[13:0], v1624[16:0], v3213[17:0]); // 3.0
    wire [24:0] v3214; shift_adder #(25, 13, 1, 1, 25, 11, 0) op_3214 (v1625[24:0], v884[12:0], v3214[24:0]); // 3.0
    wire [27:0] v3215; shift_adder #(8, 13, 1, 1, 28, -19, 0) op_3215 (v79[7:0], v884[12:0], v3215[27:0]); // 3.0
    wire [18:0] v3216; shift_adder #(11, 19, 1, 1, 19, -5, 1) op_3216 (v287[10:0], v1626[18:0], v3216[18:0]); // 3.0
    wire [18:0] v3217; shift_adder #(11, 19, 1, 1, 19, -7, 0) op_3217 (v1627[10:0], v1198[18:0], v3217[18:0]); // 3.0
    wire [13:0] v3218; shift_adder #(13, 13, 1, 1, 14, 0, 0) op_3218 (v1001[12:0], v1393[12:0], v3218[13:0]); // 3.0
    wire [19:0] v3219; shift_adder #(18, 15, 1, 1, 20, 5, 0) op_3219 (v926[17:0], v1628[14:0], v3219[19:0]); // 3.0
    wire [18:0] v3220; shift_adder #(13, 15, 1, 1, 19, -6, 1) op_3220 (v1279[12:0], v993[14:0], v3220[18:0]); // 3.0
    wire [18:0] v3221; shift_adder #(16, 15, 1, 1, 19, -3, 0) op_3221 (v1424[15:0], v1629[14:0], v3221[18:0]); // 3.0
    wire [21:0] v3222; shift_adder #(13, 15, 1, 1, 22, 7, 0) op_3222 (v1029[12:0], v1576[14:0], v3222[21:0]); // 3.0
    wire [20:0] v3223; shift_adder #(20, 16, 1, 1, 21, 4, 0) op_3223 (v1286[19:0], v1630[15:0], v3223[20:0]); // 3.0
    wire [21:0] v3224; shift_adder #(8, 12, 1, 1, 22, 10, 0) op_3224 (v120[7:0], v1631[11:0], v3224[21:0]); // 3.0
    wire [14:0] v3225; shift_adder #(13, 13, 1, 1, 15, 1, 0) op_3225 (v1324[12:0], v1202[12:0], v3225[14:0]); // 3.0
    wire [16:0] v3226; shift_adder #(11, 16, 1, 1, 17, -6, 0) op_3226 (v345[10:0], v1552[15:0], v3226[16:0]); // 3.0
    wire [23:0] v3227; shift_adder #(13, 12, 1, 1, 24, 12, 1) op_3227 (v892[12:0], v507[11:0], v3227[23:0]); // 3.0
    wire [17:0] v3228; shift_adder #(15, 13, 1, 1, 18, 5, 0) op_3228 (v1632[14:0], v1633[12:0], v3228[17:0]); // 3.0
    wire [24:0] v3229; shift_adder #(11, 25, 1, 1, 25, -11, 1) op_3229 (v413[10:0], v1634[24:0], v3229[24:0]); // 3.0
    wire [22:0] v3230; shift_adder #(21, 22, 1, 1, 23, 1, 0) op_3230 (v998[20:0], v1635[21:0], v3230[22:0]); // 3.0
    wire [16:0] v3231; shift_adder #(13, 13, 1, 1, 17, 4, 0) op_3231 (v1375[12:0], v573[12:0], v3231[16:0]); // 3.0
    wire [13:0] v3232; shift_adder #(11, 13, 1, 1, 14, -1, 0) op_3232 (v1636[10:0], v1180[12:0], v3232[13:0]); // 3.0
    wire [15:0] v3233; shift_adder #(11, 12, 1, 1, 16, 4, 1) op_3233 (v255[10:0], v1637[11:0], v3233[15:0]); // 3.0
    wire [13:0] v3234; shift_adder #(11, 13, 1, 1, 14, 1, 0) op_3234 (v1638[10:0], v1639[12:0], v3234[13:0]); // 3.0
    wire [25:0] v3235; shift_adder #(25, 12, 1, 1, 26, 14, 0) op_3235 (v829[24:0], v1640[11:0], v3235[25:0]); // 3.0
    wire [13:0] v3236; shift_adder #(12, 12, 1, 1, 14, -1, 0) op_3236 (v1641[11:0], v1642[11:0], v3236[13:0]); // 3.0
    wire [19:0] v3237; shift_adder #(13, 19, 1, 1, 20, -7, 1) op_3237 (v149[12:0], v1643[18:0], v3237[19:0]); // 3.0
    wire [18:0] v3238; shift_adder #(12, 19, 1, 1, 19, -6, 0) op_3238 (v1376[11:0], v1644[18:0], v3238[18:0]); // 3.0
    wire [36:0] v3239; shift_adder #(23, 37, 1, 1, 37, -13, 0) op_3239 (v1645[22:0], v1646[36:0], v3239[36:0]); // 3.0
    wire [28:0] v3240; shift_adder #(28, 12, 1, 1, 29, 16, 0) op_3240 (v1243[27:0], v1647[11:0], v3240[28:0]); // 3.0
    wire [24:0] v3241; shift_adder #(25, 18, 1, 1, 25, 6, 0) op_3241 (v1405[24:0], v1150[17:0], v3241[24:0]); // 3.0
    wire [24:0] v3242; shift_adder #(23, 12, 1, 1, 25, 13, 0) op_3242 (v1648[22:0], v1649[11:0], v3242[24:0]); // 3.0
    wire [18:0] v3243; shift_adder #(8, 18, 1, 1, 19, -9, 1) op_3243 (v99[7:0], v1650[17:0], v3243[18:0]); // 3.0
    wire [21:0] v3244; shift_adder #(12, 21, 1, 1, 22, -9, 0) op_3244 (v1651[11:0], v1266[20:0], v3244[21:0]); // 3.0
    wire [21:0] v3245; shift_adder #(11, 20, 1, 1, 22, 2, 1) op_3245 (v193[10:0], v1652[19:0], v3245[21:0]); // 3.0
    wire [32:0] v3246; shift_adder #(29, 32, 1, 1, 33, -3, 0) op_3246 (v1653[28:0], v1654[31:0], v3246[32:0]); // 3.0
    wire [22:0] v3247; shift_adder #(12, 22, 1, 1, 23, -10, 0) op_3247 (v1655[11:0], v1656[21:0], v3247[22:0]); // 3.0
    wire [27:0] v3248; shift_adder #(27, 12, 1, 1, 28, 15, 0) op_3248 (v1657[26:0], v1658[11:0], v3248[27:0]); // 3.0
    wire [24:0] v3249; shift_adder #(11, 12, 1, 1, 25, -14, 0) op_3249 (v270[10:0], v1659[11:0], v3249[24:0]); // 3.0
    wire [28:0] v3250; shift_adder #(12, 13, 1, 1, 29, 16, 0) op_3250 (v280[11:0], v1661[12:0], v3250[28:0]); // 3.0
    wire [25:0] v3251; shift_adder #(11, 26, 1, 1, 26, 0, 1) op_3251 (v147[10:0], v1167[25:0], v3251[25:0]); // 3.0
    wire [13:0] v3252; shift_adder #(11, 14, 1, 1, 14, -1, 1) op_3252 (v250[10:0], v1513[13:0], v3252[13:0]); // 3.0
    wire [27:0] v3253; shift_adder #(23, 27, 1, 1, 28, -4, 0) op_3253 (v1662[22:0], v1663[26:0], v3253[27:0]); // 3.0
    wire [22:0] v3254; shift_adder #(22, 13, 1, 1, 23, 9, 0) op_3254 (v1664[21:0], v1665[12:0], v3254[22:0]); // 3.0
    wire [19:0] v3255; shift_adder #(20, 11, 1, 1, 20, 5, 0) op_3255 (v1666[19:0], v941[10:0], v3255[19:0]); // 3.0
    wire [29:0] v3256; shift_adder #(9, 25, 1, 1, 30, -20, 0) op_3256 (v575[8:0], v1667[24:0], v3256[29:0]); // 3.0
    wire [22:0] v3257; shift_adder #(23, 16, 1, 1, 23, 6, 0) op_3257 (v1668[22:0], v1020[15:0], v3257[22:0]); // 3.0
    wire [12:0] v3258; shift_adder #(12, 12, 1, 1, 13, 0, 0) op_3258 (v1190[11:0], v1669[11:0], v3258[12:0]); // 3.0
    wire [15:0] v3259; shift_adder #(14, 13, 1, 1, 16, -2, 0) op_3259 (v236[13:0], v1670[12:0], v3259[15:0]); // 3.0
    wire [22:0] v3260; shift_adder #(12, 23, 1, 1, 23, -10, 0) op_3260 (v1484[11:0], v1131[22:0], v3260[22:0]); // 3.0
    wire [21:0] v3261; shift_adder #(16, 13, 1, 1, 22, -6, 1) op_3261 (v1620[15:0], v1079[12:0], v3261[21:0]); // 3.0
    wire [19:0] v3262; shift_adder #(8, 13, 1, 1, 20, -11, 1) op_3262 (v120[7:0], v1021[12:0], v3262[19:0]); // 3.0
    wire [21:0] v3263; shift_adder #(22, 17, 1, 1, 22, 3, 0) op_3263 (v1671[21:0], v1485[16:0], v3263[21:0]); // 3.0
    wire [18:0] v3264; shift_adder #(16, 14, 1, 1, 19, -3, 0) op_3264 (v1672[15:0], v1673[13:0], v3264[18:0]); // 3.0
    wire [16:0] v3265; shift_adder #(11, 17, 1, 1, 17, 0, 1) op_3265 (v175[10:0], v1674[16:0], v3265[16:0]); // 3.0
    wire [13:0] v3266; shift_adder #(11, 13, 1, 1, 14, -2, 0) op_3266 (v941[10:0], v1601[12:0], v3266[13:0]); // 3.0
    wire [17:0] v3267; shift_adder #(18, 14, 1, 1, 18, 0, 0) op_3267 (v1675[17:0], v1676[13:0], v3267[17:0]); // 3.0
    wire [14:0] v3268; shift_adder #(13, 14, 1, 1, 15, 0, 0) op_3268 (v1677[12:0], v1678[13:0], v3268[14:0]); // 3.0
    wire [15:0] v3269; shift_adder #(14, 16, 1, 1, 16, -1, 0) op_3269 (v1679[13:0], v1472[15:0], v3269[15:0]); // 3.0
    wire [20:0] v3270; shift_adder #(20, 14, 1, 1, 21, 7, 0) op_3270 (v1411[19:0], v1680[13:0], v3270[20:0]); // 3.0
    wire [18:0] v3271; shift_adder #(8, 12, 1, 1, 19, 7, 0) op_3271 (v69[7:0], v1398[11:0], v3271[18:0]); // 3.0
    wire [16:0] v3272; shift_adder #(11, 15, 1, 1, 17, -5, 0) op_3272 (v1081[10:0], v1681[14:0], v3272[16:0]); // 3.0
    wire [13:0] v3273; shift_adder #(8, 12, 1, 1, 14, -5, 1) op_3273 (v71[7:0], v1244[11:0], v3273[13:0]); // 3.0
    wire [16:0] v3274; shift_adder #(17, 16, 1, 1, 17, 0, 1) op_3274 (v887[16:0], v1682[15:0], v3274[16:0]); // 3.0
    wire [20:0] v3275; shift_adder #(20, 17, 1, 1, 21, 2, 0) op_3275 (v1683[19:0], v1684[16:0], v3275[20:0]); // 3.0
    wire [17:0] v3276; shift_adder #(11, 15, 1, 1, 18, -7, 0) op_3276 (v208[10:0], v902[14:0], v3276[17:0]); // 3.0
    wire [21:0] v3277; shift_adder #(20, 12, 1, 1, 22, 10, 0) op_3277 (v1142[19:0], v1276[11:0], v3277[21:0]); // 3.0
    wire [22:0] v3278; shift_adder #(12, 23, 1, 1, 23, -9, 0) op_3278 (v1659[11:0], v1685[22:0], v3278[22:0]); // 3.0
    wire [16:0] v3279; shift_adder #(11, 17, 1, 1, 17, -2, 0) op_3279 (v181[10:0], v1341[16:0], v3279[16:0]); // 3.0
    wire [18:0] v3280; shift_adder #(15, 17, 1, 1, 19, -3, 0) op_3280 (v1108[14:0], v1619[16:0], v3280[18:0]); // 3.0
    wire [32:0] v3281; shift_adder #(32, 12, 1, 1, 33, 20, 0) op_3281 (v1331[31:0], v1686[11:0], v3281[32:0]); // 3.0
    wire [28:0] v3282; shift_adder #(27, 15, 1, 1, 29, 13, 0) op_3282 (v1687[26:0], v1688[14:0], v3282[28:0]); // 3.0
    wire [12:0] v3283; shift_adder #(8, 12, 1, 1, 13, -3, 0) op_3283 (v101[7:0], v1689[11:0], v3283[12:0]); // 3.0
    wire [17:0] v3284; shift_adder #(15, 16, 1, 1, 18, -3, 0) op_3284 (v1690[14:0], v1691[15:0], v3284[17:0]); // 3.0
    wire [17:0] v3285; shift_adder #(8, 18, 1, 1, 18, -6, 0) op_3285 (v112[7:0], v1692[17:0], v3285[17:0]); // 3.0
    wire [31:0] v3286; shift_adder #(31, 12, 1, 1, 32, 20, 0) op_3286 (v1693[30:0], v1694[11:0], v3286[31:0]); // 3.0
    wire [19:0] v3287; shift_adder #(9, 14, 1, 1, 20, -10, 0) op_3287 (v479[8:0], v1695[13:0], v3287[19:0]); // 3.0
    wire [16:0] v3288; shift_adder #(11, 17, 1, 1, 17, -3, 1) op_3288 (v206[10:0], v972[16:0], v3288[16:0]); // 3.0
    wire [19:0] v3289; shift_adder #(11, 13, 1, 1, 20, -9, 0) op_3289 (v172[10:0], v1696[12:0], v3289[19:0]); // 3.0
    wire [19:0] v3290; shift_adder #(20, 14, 1, 1, 20, 3, 0) op_3290 (v1697[19:0], v1420[13:0], v3290[19:0]); // 3.0
    wire [27:0] v3291; shift_adder #(13, 28, 1, 1, 28, -12, 0) op_3291 (v1479[12:0], v1698[27:0], v3291[27:0]); // 3.0
    wire [19:0] v3292; shift_adder #(11, 12, 1, 1, 20, -9, 1) op_3292 (v293[10:0], v1340[11:0], v3292[19:0]); // 3.0
    wire [27:0] v3293; shift_adder #(10, 28, 1, 1, 28, -2, 1) op_3293 (v225[9:0], v1699[27:0], v3293[27:0]); // 3.0
    wire [18:0] v3294; shift_adder #(17, 19, 1, 1, 19, 0, 0) op_3294 (v1700[16:0], v1701[18:0], v3294[18:0]); // 3.0
    wire [32:0] v3295; shift_adder #(13, 13, 1, 1, 33, -20, 1) op_3295 (v920[12:0], v1189[12:0], v3295[32:0]); // 3.0
    wire [34:0] v3296; shift_adder #(34, 24, 1, 1, 35, 10, 0) op_3296 (v1702[33:0], v1703[23:0], v3296[34:0]); // 3.0
    wire [16:0] v3297; shift_adder #(13, 14, 1, 1, 17, -4, 0) op_3297 (v1704[12:0], v1705[13:0], v3297[16:0]); // 3.0
    wire [33:0] v3298; shift_adder #(13, 33, 1, 1, 34, -20, 0) op_3298 (v1706[12:0], v1707[32:0], v3298[33:0]); // 3.0
    wire [32:0] v3299; shift_adder #(10, 12, 1, 1, 33, -23, 0) op_3299 (v592[9:0], v1708[11:0], v3299[32:0]); // 3.0
    wire [28:0] v3300; shift_adder #(18, 28, 1, 1, 29, -11, 0) op_3300 (v1709[17:0], v1710[27:0], v3300[28:0]); // 3.0
    wire [14:0] v3301; shift_adder #(12, 13, 1, 1, 15, -2, 0) op_3301 (v1170[11:0], v1456[12:0], v3301[14:0]); // 3.0
    wire [11:0] v3302; shift_adder #(12, 11, 1, 1, 12, 0, 0) op_3302 (v1069[11:0], v1711[10:0], v3302[11:0]); // 3.0
    wire [35:0] v3303; shift_adder #(28, 12, 1, 1, 36, -8, 1) op_3303 (v1712[27:0], v1713[11:0], v3303[35:0]); // 3.0
    wire [22:0] v3304; shift_adder #(21, 18, 1, 1, 23, 5, 0) op_3304 (v1714[20:0], v1715[17:0], v3304[22:0]); // 3.0
    wire [15:0] v3305; shift_adder #(15, 15, 1, 1, 16, -1, 0) op_3305 (v904[14:0], v1572[14:0], v3305[15:0]); // 3.0
    wire [18:0] v3306; shift_adder #(17, 16, 1, 1, 19, -2, 0) op_3306 (v1716[16:0], v1717[15:0], v3306[18:0]); // 3.0
    wire [15:0] v3307; shift_adder #(12, 13, 1, 1, 16, -4, 1) op_3307 (v363[11:0], v985[12:0], v3307[15:0]); // 3.0
    wire [14:0] v3308; shift_adder #(11, 14, 1, 1, 15, -4, 0) op_3308 (v139[10:0], v1718[13:0], v3308[14:0]); // 3.0
    wire [15:0] v3309; shift_adder #(16, 13, 1, 1, 16, 0, 0) op_3309 (v1719[15:0], v1720[12:0], v3309[15:0]); // 3.0
    wire [21:0] v3310; shift_adder #(15, 21, 1, 1, 22, -6, 0) op_3310 (v1721[14:0], v1722[20:0], v3310[21:0]); // 3.0
    wire [31:0] v3311; shift_adder #(8, 15, 1, 1, 32, 17, 1) op_3311 (v94[7:0], v1723[14:0], v3311[31:0]); // 3.0
    wire [15:0] v3312; shift_adder #(11, 14, 1, 1, 16, 2, 0) op_3312 (v165[10:0], v1724[13:0], v3312[15:0]); // 3.0
    wire [21:0] v3313; shift_adder #(8, 15, 1, 1, 22, -13, 0) op_3313 (v118[7:0], v886[14:0], v3313[21:0]); // 3.0
    wire [27:0] v3314; shift_adder #(26, 12, 1, 1, 28, 15, 0) op_3314 (v1076[25:0], v1725[11:0], v3314[27:0]); // 3.0
    wire [28:0] v3315; shift_adder #(28, 12, 1, 1, 29, 15, 0) op_3315 (v1528[27:0], v1726[11:0], v3315[28:0]); // 3.0
    wire [30:0] v3316; shift_adder #(8, 29, 1, 1, 31, 2, 0) op_3316 (v114[7:0], v1727[28:0], v3316[30:0]); // 3.0
    wire [26:0] v3317; shift_adder #(13, 27, 1, 1, 27, -9, 0) op_3317 (v891[12:0], v1274[26:0], v3317[26:0]); // 3.0
    wire [19:0] v3318; shift_adder #(17, 17, 1, 1, 20, -3, 0) op_3318 (v1016[16:0], v917[16:0], v3318[19:0]); // 3.0
    wire [18:0] v3319; shift_adder #(19, 15, 1, 1, 19, 3, 0) op_3319 (v1643[18:0], v945[14:0], v3319[18:0]); // 3.0
    wire [22:0] v3320; shift_adder #(8, 13, 1, 1, 23, 10, 1) op_3320 (v119[7:0], v1189[12:0], v3320[22:0]); // 3.0
    wire [21:0] v3321; shift_adder #(15, 21, 1, 1, 22, -6, 0) op_3321 (v1728[14:0], v1266[20:0], v3321[21:0]); // 3.0
    wire [24:0] v3322; shift_adder #(24, 12, 1, 1, 25, 11, 0) op_3322 (v1729[23:0], v1730[11:0], v3322[24:0]); // 3.0
    wire [19:0] v3323; shift_adder #(11, 13, 1, 1, 20, 7, 1) op_3323 (v455[10:0], v1034[12:0], v3323[19:0]); // 3.0
    wire [25:0] v3324; shift_adder #(18, 25, 1, 1, 26, -7, 0) op_3324 (v1208[17:0], v1731[24:0], v3324[25:0]); // 3.0
    wire [27:0] v3325; shift_adder #(11, 25, 1, 1, 28, 3, 1) op_3325 (v341[10:0], v1732[24:0], v3325[27:0]); // 3.0
    wire [13:0] v3326; shift_adder #(8, 12, 1, 1, 14, 2, 1) op_3326 (v103[7:0], v1637[11:0], v3326[13:0]); // 3.0
    wire [22:0] v3327; shift_adder #(11, 23, 1, 1, 23, -1, 0) op_3327 (v140[10:0], v1733[22:0], v3327[22:0]); // 3.0
    wire [27:0] v3328; shift_adder #(28, 24, 1, 1, 28, 1, 0) op_3328 (v1698[27:0], v1734[23:0], v3328[27:0]); // 3.0
    wire [17:0] v3329; shift_adder #(17, 12, 1, 1, 18, 4, 0) op_3329 (v1735[16:0], v1529[11:0], v3329[17:0]); // 3.0
    wire [21:0] v3330; shift_adder #(13, 22, 1, 1, 22, -6, 0) op_3330 (v1736[12:0], v1179[21:0], v3330[21:0]); // 3.0
    wire [20:0] v3331; shift_adder #(14, 21, 1, 1, 21, -5, 0) op_3331 (v1737[13:0], v1181[20:0], v3331[20:0]); // 3.0
    wire [19:0] v3332; shift_adder #(14, 17, 1, 1, 20, -5, 0) op_3332 (v1549[13:0], v1154[16:0], v3332[19:0]); // 3.0
    wire [15:0] v3333; shift_adder #(15, 15, 1, 1, 16, 0, 0) op_3333 (v1330[14:0], v1429[14:0], v3333[15:0]); // 3.0
    wire [14:0] v3334; shift_adder #(11, 15, 1, 1, 15, -2, 0) op_3334 (v425[10:0], v1738[14:0], v3334[14:0]); // 3.0
    wire [19:0] v3335; shift_adder #(15, 20, 1, 1, 20, -1, 0) op_3335 (v1367[14:0], v1739[19:0], v3335[19:0]); // 3.0
    wire [22:0] v3336; shift_adder #(11, 15, 1, 1, 23, -12, 0) op_3336 (v156[10:0], v1740[14:0], v3336[22:0]); // 3.0
    wire [15:0] v3337; shift_adder #(11, 16, 1, 1, 16, -3, 1) op_3337 (v173[10:0], v1152[15:0], v3337[15:0]); // 3.0
    wire [19:0] v3338; shift_adder #(13, 19, 1, 1, 20, -5, 0) op_3338 (v1741[12:0], v1527[18:0], v3338[19:0]); // 3.0
    wire [22:0] v3339; shift_adder #(11, 12, 1, 1, 23, 11, 0) op_3339 (v334[10:0], v820[11:0], v3339[22:0]); // 3.0
    wire [30:0] v3340; shift_adder #(30, 11, 1, 1, 31, 19, 0) op_3340 (v984[29:0], v1742[10:0], v3340[30:0]); // 3.0
    wire [23:0] v3341; shift_adder #(12, 23, 1, 1, 24, -8, 1) op_3341 (v552[11:0], v1743[22:0], v3341[23:0]); // 3.0
    wire [23:0] v3342; shift_adder #(24, 12, 1, 1, 24, 9, 0) op_3342 (v1744[23:0], v1745[11:0], v3342[23:0]); // 3.0
    wire [29:0] v3343; shift_adder #(30, 11, 1, 1, 30, 18, 0) op_3343 (v1746[29:0], v1517[10:0], v3343[29:0]); // 3.0
    wire [21:0] v3344; shift_adder #(21, 19, 1, 1, 22, 1, 0) op_3344 (v1747[20:0], v1748[18:0], v3344[21:0]); // 3.0
    wire [14:0] v3345; shift_adder #(11, 14, 1, 1, 15, 1, 0) op_3345 (v131[10:0], v787[13:0], v3345[14:0]); // 3.0
    wire [14:0] v3346; shift_adder #(11, 14, 1, 1, 15, -2, 1) op_3346 (v246[10:0], v1749[13:0], v3346[14:0]); // 3.0
    wire [21:0] v3347; shift_adder #(18, 20, 1, 1, 22, -4, 0) op_3347 (v1750[17:0], v1101[19:0], v3347[21:0]); // 3.0
    wire [29:0] v3348; shift_adder #(12, 21, 1, 1, 30, 9, 0) op_3348 (v388[11:0], v1191[20:0], v3348[29:0]); // 3.0
    wire [25:0] v3349; shift_adder #(26, 12, 1, 1, 26, 12, 0) op_3349 (v1751[25:0], v1752[11:0], v3349[25:0]); // 3.0
    wire [24:0] v3350; shift_adder #(24, 12, 1, 1, 25, -1, 1) op_3350 (v1753[23:0], v1754[11:0], v3350[24:0]); // 3.0
    wire [21:0] v3351; shift_adder #(22, 19, 1, 1, 22, 1, 0) op_3351 (v1755[21:0], v1644[18:0], v3351[21:0]); // 3.0
    wire [19:0] v3352; shift_adder #(13, 18, 1, 1, 20, 2, 0) op_3352 (v845[12:0], v1316[17:0], v3352[19:0]); // 3.0
    wire [16:0] v3353; shift_adder #(13, 14, 1, 1, 17, -4, 1) op_3353 (v1029[12:0], v236[13:0], v3353[16:0]); // 3.0
    wire [14:0] v3354; shift_adder #(12, 15, 1, 1, 15, -1, 0) op_3354 (v1756[11:0], v1576[14:0], v3354[14:0]); // 3.0
    wire [23:0] v3355; shift_adder #(23, 13, 1, 1, 24, 10, 0) op_3355 (v1297[22:0], v1026[12:0], v3355[23:0]); // 3.0
    wire [12:0] v3356; shift_adder #(13, 12, 1, 1, 13, 0, 0) op_3356 (v920[12:0], v1370[11:0], v3356[12:0]); // 3.0
    wire [14:0] v3357; shift_adder #(12, 13, 1, 1, 15, -2, 0) op_3357 (v1757[11:0], v900[12:0], v3357[14:0]); // 3.0
    wire [14:0] v3358; shift_adder #(13, 12, 1, 1, 15, 2, 0) op_3358 (v1736[12:0], v1758[11:0], v3358[14:0]); // 3.0
    wire [23:0] v3359; shift_adder #(23, 21, 1, 1, 24, 2, 0) op_3359 (v1662[22:0], v1403[20:0], v3359[23:0]); // 3.0
    wire [22:0] v3360; shift_adder #(13, 22, 1, 1, 23, -9, 0) op_3360 (v1759[12:0], v1760[21:0], v3360[22:0]); // 3.0
    wire [17:0] v3361; shift_adder #(12, 16, 1, 1, 18, -5, 0) op_3361 (v1761[11:0], v1762[15:0], v3361[17:0]); // 3.0
    wire [32:0] v3362; shift_adder #(11, 15, 1, 1, 33, 18, 1) op_3362 (v185[10:0], v1477[14:0], v3362[32:0]); // 3.0
    wire [12:0] v3363; shift_adder #(11, 12, 1, 1, 13, 0, 1) op_3363 (v147[10:0], v1537[11:0], v3363[12:0]); // 3.0
    wire [23:0] v3364; shift_adder #(24, 14, 1, 1, 24, 5, 1) op_3364 (v1268[23:0], v603[13:0], v3364[23:0]); // 3.0
    wire [29:0] v3365; shift_adder #(30, 19, 1, 1, 30, 8, 0) op_3365 (v1763[29:0], v1764[18:0], v3365[29:0]); // 3.0
    wire [14:0] v3366; shift_adder #(14, 12, 1, 1, 15, 2, 0) op_3366 (v1281[13:0], v1765[11:0], v3366[14:0]); // 3.0
    wire [15:0] v3367; shift_adder #(14, 13, 1, 1, 16, 2, 0) op_3367 (v1380[13:0], v1766[12:0], v3367[15:0]); // 3.0
    wire [16:0] v3368; shift_adder #(13, 17, 1, 1, 17, -3, 0) op_3368 (v790[12:0], v1146[16:0], v3368[16:0]); // 3.0
    wire [13:0] v3369; shift_adder #(11, 12, 1, 1, 14, 1, 1) op_3369 (v367[10:0], v1408[11:0], v3369[13:0]); // 3.0
    wire [34:0] v3370; shift_adder #(15, 34, 1, 1, 35, -19, 0) op_3370 (v1767[14:0], v1768[33:0], v3370[34:0]); // 3.0
    wire [18:0] v3371; shift_adder #(15, 18, 1, 1, 19, -2, 0) op_3371 (v1769[14:0], v938[17:0], v3371[18:0]); // 3.0
    wire [27:0] v3372; shift_adder #(25, 28, 1, 1, 28, -2, 0) op_3372 (v1770[24:0], v1771[27:0], v3372[27:0]); // 3.0
    wire [15:0] v3373; shift_adder #(12, 14, 1, 1, 16, 2, 1) op_3373 (v434[11:0], v1104[13:0], v3373[15:0]); // 3.0
    wire [32:0] v3374; shift_adder #(19, 33, 1, 1, 33, -12, 0) op_3374 (v1772[18:0], v1773[32:0], v3374[32:0]); // 3.0
    wire [15:0] v3375; shift_adder #(15, 12, 1, 1, 16, 2, 0) op_3375 (v1774[14:0], v1775[11:0], v3375[15:0]); // 3.0
    wire [18:0] v3376; shift_adder #(11, 18, 1, 1, 19, -7, 1) op_3376 (v177[10:0], v989[17:0], v3376[18:0]); // 3.0
    wire [33:0] v3377; shift_adder #(33, 14, 1, 1, 34, 19, 0) op_3377 (v1322[32:0], v1724[13:0], v3377[33:0]); // 3.0
    wire [13:0] v3378; shift_adder #(12, 12, 1, 1, 14, 1, 0) op_3378 (v1776[11:0], v1752[11:0], v3378[13:0]); // 3.0
    wire [23:0] v3379; shift_adder #(9, 18, 1, 1, 24, -14, 0) op_3379 (v360[8:0], v1778[17:0], v3379[23:0]); // 3.0
    wire [24:0] v3380; shift_adder #(24, 14, 1, 1, 25, 10, 0) op_3380 (v1264[23:0], v976[13:0], v3380[24:0]); // 3.0
    wire [33:0] v3381; shift_adder #(33, 15, 1, 1, 34, 18, 0) op_3381 (v1779[32:0], v1780[14:0], v3381[33:0]); // 3.0
    wire [13:0] v3382; shift_adder #(12, 13, 1, 1, 14, -1, 0) op_3382 (v924[11:0], v1781[12:0], v3382[13:0]); // 3.0
    wire [17:0] v3383; shift_adder #(17, 13, 1, 1, 18, 4, 1) op_3383 (v1526[16:0], v1782[12:0], v3383[17:0]); // 3.0
    wire [14:0] v3384; shift_adder #(13, 14, 1, 1, 15, -1, 0) op_3384 (v1783[12:0], v1784[13:0], v3384[14:0]); // 3.0
    wire [36:0] v3385; shift_adder #(13, 13, 1, 1, 37, -24, 1) op_3385 (v859[12:0], v1279[12:0], v3385[36:0]); // 3.0
    wire [14:0] v3386; shift_adder #(13, 13, 1, 1, 15, -1, 0) op_3386 (v995[12:0], v813[12:0], v3386[14:0]); // 3.0
    wire [14:0] v3387; shift_adder #(11, 13, 1, 1, 15, -3, 0) op_3387 (v870[10:0], v1785[12:0], v3387[14:0]); // 3.0
    wire [19:0] v3388; shift_adder #(20, 11, 1, 1, 20, 6, 0) op_3388 (v1400[19:0], v1786[10:0], v3388[19:0]); // 3.0
    wire [14:0] v3389; shift_adder #(13, 14, 1, 1, 15, -1, 0) op_3389 (v1787[12:0], v1749[13:0], v3389[14:0]); // 3.0
    wire [20:0] v3390; shift_adder #(8, 21, 1, 1, 21, 0, 0) op_3390 (v75[7:0], v1788[20:0], v3390[20:0]); // 3.0
    wire [20:0] v3391; shift_adder #(21, 17, 1, 1, 21, 2, 0) op_3391 (v1789[20:0], v952[16:0], v3391[20:0]); // 3.0
    wire [19:0] v3392; shift_adder #(14, 19, 1, 1, 20, -6, 0) op_3392 (v1790[13:0], v547[18:0], v3392[19:0]); // 3.0
    wire [25:0] v3393; shift_adder #(13, 26, 1, 1, 26, -10, 0) op_3393 (v996[12:0], v1791[25:0], v3393[25:0]); // 3.0
    wire [20:0] v3394; shift_adder #(15, 19, 1, 1, 21, -6, 0) op_3394 (v1119[14:0], v1792[18:0], v3394[20:0]); // 3.0
    wire [13:0] v3395; shift_adder #(12, 12, 1, 1, 14, -1, 0) op_3395 (v1262[11:0], v1025[11:0], v3395[13:0]); // 3.0
    wire [15:0] v3396; shift_adder #(15, 9, 1, 1, 16, 5, 1) op_3396 (v1015[14:0], v479[8:0], v3396[15:0]); // 3.0
    wire [16:0] v3397; shift_adder #(11, 17, 1, 1, 17, -1, 0) op_3397 (v266[10:0], v876[16:0], v3397[16:0]); // 3.0
    wire [16:0] v3398; shift_adder #(16, 14, 1, 1, 17, 2, 0) op_3398 (v1793[15:0], v1794[13:0], v3398[16:0]); // 3.0
    wire [15:0] v3399; shift_adder #(13, 16, 1, 1, 16, 0, 0) op_3399 (v1393[12:0], v1795[15:0], v3399[15:0]); // 3.0
    wire [22:0] v3400; shift_adder #(13, 23, 1, 1, 23, -6, 0) op_3400 (v1796[12:0], v1797[22:0], v3400[22:0]); // 3.0
    wire [23:0] v3401; shift_adder #(23, 13, 1, 1, 24, 11, 0) op_3401 (v1798[22:0], v1799[12:0], v3401[23:0]); // 3.0
    wire [18:0] v3402; shift_adder #(8, 11, 1, 1, 19, 8, 0) op_3402 (v76[7:0], v1800[10:0], v3402[18:0]); // 3.0
    wire [20:0] v3403; shift_adder #(16, 19, 1, 1, 21, 2, 0) op_3403 (v504[15:0], v1643[18:0], v3403[20:0]); // 3.0
    wire [18:0] v3404; shift_adder #(12, 19, 1, 1, 19, -1, 0) op_3404 (v385[11:0], v1801[18:0], v3404[18:0]); // 3.0
    wire [15:0] v3405; shift_adder #(12, 12, 1, 1, 16, 4, 0) op_3405 (v257[11:0], v1262[11:0], v3405[15:0]); // 3.0
    wire [17:0] v3406; shift_adder #(9, 12, 1, 1, 18, -8, 0) op_3406 (v395[8:0], v1589[11:0], v3406[17:0]); // 3.0
    wire [16:0] v3407; shift_adder #(15, 13, 1, 1, 17, 3, 0) op_3407 (v1767[14:0], v1802[12:0], v3407[16:0]); // 3.0
    wire [29:0] v3408; shift_adder #(28, 23, 1, 1, 30, 6, 0) op_3408 (v1803[27:0], v980[22:0], v3408[29:0]); // 3.0
    wire [26:0] v3409; shift_adder #(15, 27, 1, 1, 27, -10, 0) op_3409 (v905[14:0], v1246[26:0], v3409[26:0]); // 3.0
    wire [19:0] v3410; shift_adder #(11, 13, 1, 1, 20, -9, 0) op_3410 (v317[10:0], v1180[12:0], v3410[19:0]); // 3.0
    wire [17:0] v3411; shift_adder #(15, 17, 1, 1, 18, -1, 0) op_3411 (v840[14:0], v1804[16:0], v3411[17:0]); // 3.0
    wire [20:0] v3412; shift_adder #(19, 12, 1, 1, 21, 8, 0) op_3412 (v1805[18:0], v1806[11:0], v3412[20:0]); // 3.0
    wire [18:0] v3413; shift_adder #(11, 13, 1, 1, 19, 6, 1) op_3413 (v259[10:0], v1134[12:0], v3413[18:0]); // 3.0
    wire [24:0] v3414; shift_adder #(8, 24, 1, 1, 25, -16, 1) op_3414 (v81[7:0], v1807[23:0], v3414[24:0]); // 3.0
    wire [27:0] v3415; shift_adder #(11, 24, 1, 1, 28, 4, 1) op_3415 (v233[10:0], v1808[23:0], v3415[27:0]); // 3.0
    wire [18:0] v3416; shift_adder #(17, 17, 1, 1, 19, 2, 0) op_3416 (v1809[16:0], v1455[16:0], v3416[18:0]); // 3.0
    wire [11:0] v3417; shift_adder #(8, 11, 1, 1, 12, -2, 1) op_3417 (v73[7:0], v1810[10:0], v3417[11:0]); // 3.0
    wire [35:0] v3418; shift_adder #(14, 11, 1, 1, 36, 25, 1) op_3418 (v1165[13:0], v213[10:0], v3418[35:0]); // 3.0
    wire [14:0] v3419; shift_adder #(13, 13, 1, 1, 15, 2, 0) op_3419 (v1202[12:0], v1811[12:0], v3419[14:0]); // 3.0
    wire [15:0] v3420; shift_adder #(15, 15, 1, 1, 16, 1, 0) op_3420 (v1812[14:0], v1124[14:0], v3420[15:0]); // 3.0
    wire [12:0] v3421; shift_adder #(11, 11, 1, 1, 13, -2, 1) op_3421 (v323[10:0], v1284[10:0], v3421[12:0]); // 3.0
    wire [18:0] v3422; shift_adder #(14, 19, 1, 1, 19, -4, 0) op_3422 (v1813[13:0], v1814[18:0], v3422[18:0]); // 3.0
    wire [32:0] v3423; shift_adder #(17, 32, 1, 1, 33, -16, 0) op_3423 (v1716[16:0], v1815[31:0], v3423[32:0]); // 3.0
    wire [21:0] v3424; shift_adder #(22, 16, 1, 1, 22, 5, 0) op_3424 (v918[21:0], v1816[15:0], v3424[21:0]); // 3.0
    wire [18:0] v3425; shift_adder #(14, 19, 1, 1, 19, -4, 0) op_3425 (v1817[13:0], v1530[18:0], v3425[18:0]); // 3.0
    wire [28:0] v3426; shift_adder #(14, 28, 1, 1, 29, -14, 0) op_3426 (v1818[13:0], v1710[27:0], v3426[28:0]); // 3.0
    wire [17:0] v3427; shift_adder #(13, 18, 1, 1, 18, -4, 0) op_3427 (v1819[12:0], v1820[17:0], v3427[17:0]); // 3.0
    wire [13:0] v3428; shift_adder #(12, 12, 1, 1, 14, -2, 0) op_3428 (v1821[11:0], v1822[11:0], v3428[13:0]); // 3.0
    wire [22:0] v3429; shift_adder #(21, 20, 1, 1, 23, -1, 0) op_3429 (v1823[20:0], v1824[19:0], v3429[22:0]); // 3.0
    wire [14:0] v3430; shift_adder #(13, 13, 1, 1, 15, -2, 0) op_3430 (v920[12:0], v1825[12:0], v3430[14:0]); // 3.0
    wire [22:0] v3431; shift_adder #(11, 19, 1, 1, 23, -12, 1) op_3431 (v374[10:0], v1826[18:0], v3431[22:0]); // 3.0
    wire [16:0] v3432; shift_adder #(10, 16, 1, 1, 17, 1, 0) op_3432 (v501[9:0], v1827[15:0], v3432[16:0]); // 3.0
    wire [14:0] v3433; shift_adder #(15, 12, 1, 1, 15, 1, 0) op_3433 (v1828[14:0], v1829[11:0], v3433[14:0]); // 3.0
    wire [19:0] v3434; shift_adder #(19, 19, 1, 1, 20, 0, 0) op_3434 (v1036[18:0], v1830[18:0], v3434[19:0]); // 3.0
    wire [17:0] v3435; shift_adder #(12, 16, 1, 1, 18, -5, 0) op_3435 (v1399[11:0], v1831[15:0], v3435[17:0]); // 3.0
    wire [15:0] v3436; shift_adder #(13, 15, 1, 1, 16, -2, 0) op_3436 (v1177[12:0], v1430[14:0], v3436[15:0]); // 3.0
    wire [15:0] v3437; shift_adder #(11, 10, 1, 1, 16, 6, 0) op_3437 (v772[10:0], v254[9:0], v3437[15:0]); // 3.0
    wire [15:0] v3438; shift_adder #(11, 15, 1, 1, 16, -5, 0) op_3438 (v358[10:0], v1832[14:0], v3438[15:0]); // 3.0
    wire [15:0] v3439; shift_adder #(15, 14, 1, 1, 16, 1, 0) op_3439 (v1833[14:0], v1834[13:0], v3439[15:0]); // 3.0
    wire [14:0] v3440; shift_adder #(13, 12, 1, 1, 15, -2, 0) op_3440 (v1349[12:0], v808[11:0], v3440[14:0]); // 3.0
    wire [23:0] v3441; shift_adder #(24, 18, 1, 1, 24, 5, 0) op_3441 (v1058[23:0], v1835[17:0], v3441[23:0]); // 3.0
    wire [14:0] v3442; shift_adder #(12, 14, 1, 1, 15, -2, 0) op_3442 (v1836[11:0], v1135[13:0], v3442[14:0]); // 3.0
    wire [14:0] v3443; shift_adder #(11, 14, 1, 1, 15, 1, 0) op_3443 (v173[10:0], v964[13:0], v3443[14:0]); // 3.0
    wire [25:0] v3444; shift_adder #(12, 24, 1, 1, 26, -13, 0) op_3444 (v1234[11:0], v1837[23:0], v3444[25:0]); // 3.0
    wire [15:0] v3445; shift_adder #(12, 15, 1, 1, 16, -4, 0) op_3445 (v1043[11:0], v781[14:0], v3445[15:0]); // 3.0
    wire [15:0] v3446; shift_adder #(12, 15, 1, 1, 16, -3, 0) op_3446 (v1262[11:0], v904[14:0], v3446[15:0]); // 3.0
    wire [25:0] v3447; shift_adder #(8, 26, 1, 1, 26, -8, 1) op_3447 (v85[7:0], v1838[25:0], v3447[25:0]); // 3.0
    wire [19:0] v3448; shift_adder #(11, 13, 1, 1, 20, 7, 0) op_3448 (v275[10:0], v813[12:0], v3448[19:0]); // 3.0
    wire [21:0] v3449; shift_adder #(11, 14, 1, 1, 22, 8, 0) op_3449 (v142[10:0], v830[13:0], v3449[21:0]); // 3.0
    wire [23:0] v3450; shift_adder #(12, 24, 1, 1, 24, -5, 0) op_3450 (v409[11:0], v1839[23:0], v3450[23:0]); // 3.0
    wire [23:0] v3451; shift_adder #(21, 23, 1, 1, 24, -3, 0) op_3451 (v1062[20:0], v1733[22:0], v3451[23:0]); // 3.0
    wire [15:0] v3452; shift_adder #(16, 13, 1, 1, 16, 1, 0) op_3452 (v1840[15:0], v1421[12:0], v3452[15:0]); // 3.0
    wire [25:0] v3453; shift_adder #(25, 13, 1, 1, 26, 12, 0) op_3453 (v1444[24:0], v795[12:0], v3453[25:0]); // 3.0
    wire [24:0] v3454; shift_adder #(17, 24, 1, 1, 25, -7, 0) op_3454 (v887[16:0], v1753[23:0], v3454[24:0]); // 3.0
    wire [17:0] v3455; shift_adder #(18, 14, 1, 1, 18, 3, 0) op_3455 (v1841[17:0], v1135[13:0], v3455[17:0]); // 3.0
    wire [24:0] v3456; shift_adder #(23, 22, 1, 1, 25, 2, 0) op_3456 (v1842[22:0], v1843[21:0], v3456[24:0]); // 3.0
    wire [24:0] v3457; shift_adder #(9, 19, 1, 1, 25, -15, 1) op_3457 (v256[8:0], v1764[18:0], v3457[24:0]); // 3.0
    wire [18:0] v3458; shift_adder #(8, 15, 1, 1, 19, -10, 1) op_3458 (v77[7:0], v779[14:0], v3458[18:0]); // 3.0
    wire [13:0] v3459; shift_adder #(11, 13, 1, 1, 14, -1, 1) op_3459 (v185[10:0], v1551[12:0], v3459[13:0]); // 3.0
    wire [20:0] v3460; shift_adder #(17, 20, 1, 1, 21, -3, 0) op_3460 (v1146[16:0], v1844[19:0], v3460[20:0]); // 3.0
    wire [25:0] v3461; shift_adder #(26, 18, 1, 1, 26, 5, 0) op_3461 (v1845[25:0], v1846[17:0], v3461[25:0]); // 3.0
    wire [17:0] v3462; shift_adder #(14, 17, 1, 1, 18, -2, 0) op_3462 (v1072[13:0], v1847[16:0], v3462[17:0]); // 3.0
    wire [18:0] v3463; shift_adder #(15, 12, 1, 1, 19, 7, 0) op_3463 (v1583[14:0], v1398[11:0], v3463[18:0]); // 3.0
    wire [17:0] v3464; shift_adder #(12, 11, 1, 1, 18, -6, 1) op_3464 (v183[11:0], v1161[10:0], v3464[17:0]); // 3.0
    wire [19:0] v3465; shift_adder #(11, 19, 1, 1, 20, -8, 1) op_3465 (v219[10:0], v1848[18:0], v3465[19:0]); // 3.0
    wire [18:0] v3466; shift_adder #(17, 15, 1, 1, 19, 4, 0) op_3466 (v1392[16:0], v1849[14:0], v3466[18:0]); // 3.0
    wire [16:0] v3467; shift_adder #(15, 12, 1, 1, 17, 4, 0) op_3467 (v1120[14:0], v1850[11:0], v3467[16:0]); // 3.0
    wire [25:0] v3468; shift_adder #(26, 17, 1, 1, 26, 7, 0) op_3468 (v1845[25:0], v832[16:0], v3468[25:0]); // 3.0
    wire [19:0] v3469; shift_adder #(18, 12, 1, 1, 20, 7, 0) op_3469 (v1851[17:0], v1852[11:0], v3469[19:0]); // 3.0
    wire [18:0] v3470; shift_adder #(8, 13, 1, 1, 19, 6, 0) op_3470 (v65[7:0], v1853[12:0], v3470[18:0]); // 3.0
    wire [16:0] v3471; shift_adder #(11, 17, 1, 1, 17, -1, 0) op_3471 (v785[10:0], v1542[16:0], v3471[16:0]); // 3.0
    wire [27:0] v3472; shift_adder #(27, 17, 1, 1, 28, 11, 0) op_3472 (v1854[26:0], v1151[16:0], v3472[27:0]); // 3.0
    wire [25:0] v3473; shift_adder #(18, 25, 1, 1, 26, -7, 0) op_3473 (v1391[17:0], v916[24:0], v3473[25:0]); // 3.0
    wire [26:0] v3474; shift_adder #(11, 13, 1, 1, 27, 14, 0) op_3474 (v303[10:0], v833[12:0], v3474[26:0]); // 3.0
    wire [21:0] v3475; shift_adder #(13, 22, 1, 1, 22, -8, 0) op_3475 (v1508[12:0], v1855[21:0], v3475[21:0]); // 3.0
    wire [23:0] v3476; shift_adder #(12, 23, 1, 1, 24, -10, 0) op_3476 (v1856[11:0], v1857[22:0], v3476[23:0]); // 3.0
    wire [18:0] v3477; shift_adder #(15, 18, 1, 1, 19, -4, 0) op_3477 (v1858[14:0], v1841[17:0], v3477[18:0]); // 3.0
    wire [19:0] v3478; shift_adder #(14, 20, 1, 1, 20, -4, 0) op_3478 (v1859[13:0], v1860[19:0], v3478[19:0]); // 3.0
    wire [21:0] v3479; shift_adder #(11, 12, 1, 1, 22, -11, 1) op_3479 (v1049[10:0], v1862[11:0], v3479[21:0]); // 3.0
    wire [13:0] v3480; shift_adder #(13, 12, 1, 1, 14, 1, 0) op_3480 (v1863[12:0], v1566[11:0], v3480[13:0]); // 3.0
    wire [27:0] v3481; shift_adder #(8, 21, 1, 1, 28, 7, 1) op_3481 (v103[7:0], v1864[20:0], v3481[27:0]); // 3.0
    wire [13:0] v3482; shift_adder #(13, 12, 1, 1, 14, 0, 0) op_3482 (v1385[12:0], v1865[11:0], v3482[13:0]); // 3.0
    wire [17:0] v3483; shift_adder #(8, 12, 1, 1, 18, -9, 1) op_3483 (v66[7:0], v1866[11:0], v3483[17:0]); // 3.0
    wire [15:0] v3484; shift_adder #(15, 14, 1, 1, 16, 1, 0) op_3484 (v1867[14:0], v1162[13:0], v3484[15:0]); // 3.0
    wire [15:0] v3485; shift_adder #(15, 15, 1, 1, 16, 0, 0) op_3485 (v1477[14:0], v1429[14:0], v3485[15:0]); // 3.0
    wire [17:0] v3486; shift_adder #(17, 12, 1, 1, 18, 6, 0) op_3486 (v1618[16:0], v1031[11:0], v3486[17:0]); // 3.0
    wire [19:0] v3487; shift_adder #(11, 13, 1, 1, 20, -9, 0) op_3487 (v229[10:0], v793[12:0], v3487[19:0]); // 3.0
    wire [16:0] v3488; shift_adder #(16, 15, 1, 1, 17, -1, 0) op_3488 (v1795[15:0], v1252[14:0], v3488[16:0]); // 3.0
    wire [17:0] v3489; shift_adder #(9, 13, 1, 1, 18, -8, 0) op_3489 (v360[8:0], v1500[12:0], v3489[17:0]); // 3.0
    wire [18:0] v3490; shift_adder #(11, 18, 1, 1, 19, -7, 0) op_3490 (v1868[10:0], v1869[17:0], v3490[18:0]); // 3.0
    wire [33:0] v3491; shift_adder #(21, 34, 1, 1, 34, -11, 0) op_3491 (v1062[20:0], v1870[33:0], v3491[33:0]); // 3.0
    wire [33:0] v3492; shift_adder #(12, 10, 1, 1, 34, -22, 1) op_3492 (v1571[11:0], v632[9:0], v3492[33:0]); // 3.0
    wire [32:0] v3493; shift_adder #(12, 12, 1, 1, 33, -21, 1) op_3493 (v1399[11:0], v1871[11:0], v3493[32:0]); // 3.0
    wire [36:0] v3494; shift_adder #(13, 12, 1, 1, 37, 25, 1) op_3494 (v1021[12:0], v402[11:0], v3494[36:0]); // 3.0
    wire [15:0] v3495; shift_adder #(11, 13, 1, 1, 16, -5, 0) op_3495 (v361[10:0], v1872[12:0], v3495[15:0]); // 3.0
    wire [13:0] v3496; shift_adder #(12, 12, 1, 1, 14, -1, 0) op_3496 (v1873[11:0], v965[11:0], v3496[13:0]); // 3.0
    wire [15:0] v3497; shift_adder #(15, 14, 1, 1, 16, 1, 0) op_3497 (v1874[14:0], v1112[13:0], v3497[15:0]); // 3.0
    wire [32:0] v3498; shift_adder #(25, 33, 1, 1, 33, -7, 0) op_3498 (v1875[24:0], v1876[32:0], v3498[32:0]); // 3.0
    wire [12:0] v3499; shift_adder #(12, 11, 1, 1, 13, 0, 0) op_3499 (v1462[11:0], v1877[10:0], v3499[12:0]); // 3.0
    wire [13:0] v3500; shift_adder #(13, 13, 1, 1, 14, 0, 0) op_3500 (v1479[12:0], v995[12:0], v3500[13:0]); // 3.0
    wire [21:0] v3501; shift_adder #(16, 22, 1, 1, 22, -1, 1) op_3501 (v1213[15:0], v587[21:0], v3501[21:0]); // 3.0
    wire [21:0] v3502; shift_adder #(21, 13, 1, 1, 22, 8, 0) op_3502 (v1144[20:0], v1825[12:0], v3502[21:0]); // 3.0
    wire [26:0] v3503; shift_adder #(8, 27, 1, 1, 27, -7, 0) op_3503 (v111[7:0], v1878[26:0], v3503[26:0]); // 3.0
    wire [29:0] v3504; shift_adder #(30, 15, 1, 1, 30, 14, 0) op_3504 (v1746[29:0], v1879[14:0], v3504[29:0]); // 3.0
    wire [12:0] v3505; shift_adder #(12, 12, 1, 1, 13, 0, 0) op_3505 (v1211[11:0], v835[11:0], v3505[12:0]); // 3.0
    wire [25:0] v3506; shift_adder #(8, 14, 1, 1, 26, -17, 0) op_3506 (v111[7:0], v1135[13:0], v3506[25:0]); // 3.0
    wire [15:0] v3507; shift_adder #(12, 15, 1, 1, 16, -4, 0) op_3507 (v1031[11:0], v1880[14:0], v3507[15:0]); // 3.0
    wire [21:0] v3508; shift_adder #(11, 12, 1, 1, 22, 10, 1) op_3508 (v242[10:0], v1686[11:0], v3508[21:0]); // 3.0
    wire [26:0] v3509; shift_adder #(12, 26, 1, 1, 27, -14, 0) op_3509 (v1570[11:0], v1881[25:0], v3509[26:0]); // 3.0
    wire [23:0] v3510; shift_adder #(17, 18, 1, 1, 24, -7, 0) op_3510 (v1175[16:0], v989[17:0], v3510[23:0]); // 3.0
    wire [25:0] v3511; shift_adder #(12, 13, 1, 1, 26, 13, 0) op_3511 (v397[11:0], v1280[12:0], v3511[25:0]); // 3.0
    wire [28:0] v3512; shift_adder #(21, 26, 1, 1, 29, -8, 0) op_3512 (v1181[20:0], v1882[25:0], v3512[28:0]); // 3.0
    wire [19:0] v3513; shift_adder #(17, 18, 1, 1, 20, 2, 0) op_3513 (v1883[16:0], v1715[17:0], v3513[19:0]); // 3.0
    wire [17:0] v3514; shift_adder #(18, 13, 1, 1, 18, 2, 0) op_3514 (v1884[17:0], v1407[12:0], v3514[17:0]); // 3.0
    wire [13:0] v3515; shift_adder #(9, 13, 1, 1, 14, -4, 1) op_3515 (v309[8:0], v1346[12:0], v3515[13:0]); // 3.0
    wire [21:0] v3516; shift_adder #(8, 22, 1, 1, 22, -10, 1) op_3516 (v106[7:0], v1885[21:0], v3516[21:0]); // 3.0
    wire [24:0] v3517; shift_adder #(8, 20, 1, 1, 25, 5, 1) op_3517 (v65[7:0], v1886[19:0], v3517[24:0]); // 3.0
    wire [22:0] v3518; shift_adder #(16, 18, 1, 1, 23, -7, 0) op_3518 (v1887[15:0], v1445[17:0], v3518[22:0]); // 3.0
    wire [16:0] v3519; shift_adder #(12, 12, 1, 1, 17, -5, 0) op_3519 (v1309[11:0], v1888[11:0], v3519[16:0]); // 3.0
    wire [18:0] v3520; shift_adder #(16, 18, 1, 1, 19, -2, 0) op_3520 (v1889[15:0], v1890[17:0], v3520[18:0]); // 3.0
    wire [15:0] v3521; shift_adder #(14, 13, 1, 1, 16, 2, 0) op_3521 (v1891[13:0], v1892[12:0], v3521[15:0]); // 3.0
    wire [20:0] v3522; shift_adder #(8, 12, 1, 1, 21, 9, 1) op_3522 (v69[7:0], v1893[11:0], v3522[20:0]); // 3.0
    wire [17:0] v3523; shift_adder #(9, 18, 1, 1, 18, -5, 1) op_3523 (v486[8:0], v1890[17:0], v3523[17:0]); // 3.0
    wire [12:0] v3524; shift_adder #(11, 13, 1, 1, 13, 0, 1) op_3524 (v269[10:0], v1560[12:0], v3524[12:0]); // 3.0
    wire [21:0] v3525; shift_adder #(17, 11, 1, 1, 22, 10, 0) op_3525 (v1037[16:0], v1894[10:0], v3525[21:0]); // 3.0
    wire [21:0] v3526; shift_adder #(18, 21, 1, 1, 22, -3, 1) op_3526 (v968[17:0], v1895[20:0], v3526[21:0]); // 3.0
    wire [13:0] v3527; shift_adder #(13, 12, 1, 1, 14, 1, 0) op_3527 (v1375[12:0], v1125[11:0], v3527[13:0]); // 3.0
    wire [32:0] v3528; shift_adder #(32, 16, 1, 1, 33, 16, 0) op_3528 (v1896[31:0], v1897[15:0], v3528[32:0]); // 3.0
    wire [16:0] v3529; shift_adder #(12, 16, 1, 1, 17, -3, 0) op_3529 (v1898[11:0], v1899[15:0], v3529[16:0]); // 3.0
    wire [21:0] v3530; shift_adder #(11, 15, 1, 1, 22, 7, 1) op_3530 (v353[10:0], v1812[14:0], v3530[21:0]); // 3.0
    wire [19:0] v3531; shift_adder #(19, 13, 1, 1, 20, 6, 0) op_3531 (v1900[18:0], v1901[12:0], v3531[19:0]); // 3.0
    wire [19:0] v3532; shift_adder #(8, 20, 1, 1, 20, -9, 0) op_3532 (v91[7:0], v1902[19:0], v3532[19:0]); // 3.0
    wire [32:0] v3533; shift_adder #(30, 26, 1, 1, 33, 7, 0) op_3533 (v1223[29:0], v1791[25:0], v3533[32:0]); // 3.0
    wire [22:0] v3534; shift_adder #(13, 14, 1, 1, 23, 9, 0) op_3534 (v344[12:0], v1749[13:0], v3534[22:0]); // 3.0
    wire [18:0] v3535; shift_adder #(13, 18, 1, 1, 19, -5, 0) op_3535 (v845[12:0], v939[17:0], v3535[18:0]); // 3.0
    wire [23:0] v3536; shift_adder #(23, 13, 1, 1, 24, 9, 0) op_3536 (v1903[22:0], v795[12:0], v3536[23:0]); // 3.0
    wire [37:0] v3537; shift_adder #(15, 11, 1, 1, 38, 27, 1) op_3537 (v1904[14:0], v636[10:0], v3537[37:0]); // 3.0
    wire [19:0] v3538; shift_adder #(18, 11, 1, 1, 20, 8, 0) op_3538 (v1451[17:0], v1905[10:0], v3538[19:0]); // 3.0
    wire [39:0] v3539; shift_adder #(12, 13, 1, 1, 40, -28, 1) op_3539 (v1906[11:0], v1907[12:0], v3539[39:0]); // 3.0
    wire [15:0] v3540; shift_adder #(13, 13, 1, 1, 16, 2, 0) op_3540 (v1908[12:0], v1909[12:0], v3540[15:0]); // 3.0
    wire [18:0] v3541; shift_adder #(12, 17, 1, 1, 19, -6, 0) op_3541 (v801[11:0], v1910[16:0], v3541[18:0]); // 3.0
    wire [12:0] v3542; shift_adder #(8, 13, 1, 1, 13, -1, 0) op_3542 (v111[7:0], v1741[12:0], v3542[12:0]); // 3.0
    wire [17:0] v3543; shift_adder #(13, 16, 1, 1, 18, -4, 0) op_3543 (v1911[12:0], v1912[15:0], v3543[17:0]); // 3.0
    wire [16:0] v3544; shift_adder #(16, 13, 1, 1, 17, 2, 0) op_3544 (v1913[15:0], v1914[12:0], v3544[16:0]); // 3.0
    wire [16:0] v3545; shift_adder #(17, 13, 1, 1, 17, 2, 0) op_3545 (v1674[16:0], v915[12:0], v3545[16:0]); // 3.0
    wire [15:0] v3546; shift_adder #(12, 13, 1, 1, 16, 3, 0) op_3546 (v174[11:0], v1295[12:0], v3546[15:0]); // 3.0
    wire [13:0] v3547; shift_adder #(12, 13, 1, 1, 14, 0, 0) op_3547 (v1915[11:0], v1326[12:0], v3547[13:0]); // 3.0
    wire [13:0] v3548; shift_adder #(12, 12, 1, 1, 14, -1, 0) op_3548 (v1888[11:0], v1537[11:0], v3548[13:0]); // 3.0
    wire [15:0] v3549; shift_adder #(15, 13, 1, 1, 16, 3, 0) op_3549 (v922[14:0], v1916[12:0], v3549[15:0]); // 3.0
    wire [17:0] v3550; shift_adder #(17, 13, 1, 1, 18, 4, 0) op_3550 (v1684[16:0], v1422[12:0], v3550[17:0]); // 3.0
    wire [35:0] v3551; shift_adder #(19, 34, 1, 1, 36, -16, 0) op_3551 (v1917[18:0], v1918[33:0], v3551[35:0]); // 3.0
    wire [20:0] v3552; shift_adder #(21, 15, 1, 1, 21, 2, 1) op_3552 (v951[20:0], v1919[14:0], v3552[20:0]); // 3.0
    wire [20:0] v3553; shift_adder #(20, 18, 1, 1, 21, 2, 0) op_3553 (v1224[19:0], v1094[17:0], v3553[20:0]); // 3.0
    wire [19:0] v3554; shift_adder #(15, 19, 1, 1, 20, -5, 1) op_3554 (v993[14:0], v1848[18:0], v3554[19:0]); // 3.0
    wire [15:0] v3555; shift_adder #(16, 12, 1, 1, 16, 1, 0) op_3555 (v1920[15:0], v873[11:0], v3555[15:0]); // 3.0
    wire [14:0] v3556; shift_adder #(15, 12, 1, 1, 15, 1, 0) op_3556 (v1921[14:0], v1922[11:0], v3556[14:0]); // 3.0
    wire [13:0] v3557; shift_adder #(10, 12, 1, 1, 14, 2, 0) op_3557 (v366[9:0], v1923[11:0], v3557[13:0]); // 3.0
    wire [30:0] v3558; shift_adder #(17, 13, 1, 1, 31, 18, 1) op_3558 (v1063[16:0], v1924[12:0], v3558[30:0]); // 3.0
    wire [27:0] v3559; shift_adder #(10, 25, 1, 1, 28, 3, 0) op_3559 (v461[9:0], v1925[24:0], v3559[27:0]); // 3.0
    wire [31:0] v3560; shift_adder #(8, 11, 1, 1, 32, -23, 1) op_3560 (v123[7:0], v1395[10:0], v3560[31:0]); // 3.0
    wire [21:0] v3561; shift_adder #(21, 14, 1, 1, 22, 7, 0) op_3561 (v1926[20:0], v1927[13:0], v3561[21:0]); // 3.0
    wire [17:0] v3562; shift_adder #(16, 16, 1, 1, 18, -1, 0) op_3562 (v1928[15:0], v1929[15:0], v3562[17:0]); // 3.0
    wire [27:0] v3563; shift_adder #(11, 23, 1, 1, 28, 5, 0) op_3563 (v319[10:0], v1141[22:0], v3563[27:0]); // 3.0
    wire [27:0] v3564; shift_adder #(17, 23, 1, 1, 28, -11, 1) op_3564 (v1151[16:0], v1930[22:0], v3564[27:0]); // 3.0
    wire [27:0] v3565; shift_adder #(21, 25, 1, 1, 28, -7, 0) op_3565 (v1090[20:0], v1634[24:0], v3565[27:0]); // 3.0
    wire [20:0] v3566; shift_adder #(13, 16, 1, 1, 21, 5, 0) op_3566 (v149[12:0], v1425[15:0], v3566[20:0]); // 3.0
    wire [31:0] v3567; shift_adder #(13, 11, 1, 1, 32, 21, 1) op_3567 (v882[12:0], v644[10:0], v3567[31:0]); // 3.0
    wire [23:0] v3568; shift_adder #(19, 22, 1, 1, 24, -5, 0) op_3568 (v1931[18:0], v1388[21:0], v3568[23:0]); // 3.0
    wire [16:0] v3569; shift_adder #(13, 15, 1, 1, 17, 2, 0) op_3569 (v344[12:0], v1932[14:0], v3569[16:0]); // 3.0
    wire [24:0] v3570; shift_adder #(11, 17, 1, 1, 25, -14, 0) op_3570 (v234[10:0], v1467[16:0], v3570[24:0]); // 3.0
    wire [14:0] v3571; shift_adder #(15, 14, 1, 1, 15, 0, 0) op_3571 (v1933[14:0], v842[13:0], v3571[14:0]); // 3.0
    wire [15:0] v3572; shift_adder #(14, 11, 1, 1, 16, 4, 0) op_3572 (v1934[13:0], v1419[10:0], v3572[15:0]); // 3.0
    wire [19:0] v3573; shift_adder #(20, 18, 1, 1, 20, 1, 0) op_3573 (v1224[19:0], v1561[17:0], v3573[19:0]); // 3.0
    wire [17:0] v3574; shift_adder #(14, 16, 1, 1, 18, -3, 0) op_3574 (v1290[13:0], v1249[15:0], v3574[17:0]); // 3.0
    wire [26:0] v3575; shift_adder #(15, 25, 1, 1, 27, -12, 0) op_3575 (v922[14:0], v1935[24:0], v3575[26:0]); // 3.0
    wire [19:0] v3576; shift_adder #(14, 12, 1, 1, 20, 8, 1) op_3576 (v249[13:0], v1558[11:0], v3576[19:0]); // 3.0
    wire [15:0] v3577; shift_adder #(12, 12, 1, 1, 16, 4, 1) op_3577 (v867[11:0], v824[11:0], v3577[15:0]); // 3.0
    wire [25:0] v3578; shift_adder #(22, 19, 1, 1, 26, 7, 0) op_3578 (v1342[21:0], v1195[18:0], v3578[25:0]); // 3.0
    wire [28:0] v3579; shift_adder #(14, 9, 1, 1, 29, -15, 0) op_3579 (v1695[13:0], v384[8:0], v3579[28:0]); // 3.0
    wire [23:0] v3580; shift_adder #(23, 12, 1, 1, 24, 10, 0) op_3580 (v1936[22:0], v1537[11:0], v3580[23:0]); // 3.0
    wire [28:0] v3581; shift_adder #(14, 28, 1, 1, 29, -14, 0) op_3581 (v1139[13:0], v1245[27:0], v3581[28:0]); // 3.0
    wire [14:0] v3582; shift_adder #(11, 15, 1, 1, 15, -3, 0) op_3582 (v182[10:0], v1681[14:0], v3582[14:0]); // 3.0
    wire [24:0] v3583; shift_adder #(8, 15, 1, 1, 25, 10, 1) op_3583 (v124[7:0], v1774[14:0], v3583[24:0]); // 3.0
    wire [13:0] v3584; shift_adder #(13, 13, 1, 1, 14, 0, 0) op_3584 (v1482[12:0], v834[12:0], v3584[13:0]); // 3.0
    wire [16:0] v3585; shift_adder #(13, 17, 1, 1, 17, -3, 1) op_3585 (v826[12:0], v1937[16:0], v3585[16:0]); // 3.0
    wire [18:0] v3586; shift_adder #(18, 14, 1, 1, 19, 4, 0) op_3586 (v1938[17:0], v1939[13:0], v3586[18:0]); // 3.0
    wire [14:0] v3587; shift_adder #(14, 12, 1, 1, 15, 2, 0) op_3587 (v1014[13:0], v1940[11:0], v3587[14:0]); // 3.0
    wire [14:0] v3588; shift_adder #(15, 13, 1, 1, 15, 0, 0) op_3588 (v1576[14:0], v1941[12:0], v3588[14:0]); // 3.0
    wire [20:0] v3589; shift_adder #(21, 19, 1, 1, 21, 0, 0) op_3589 (v1090[20:0], v1942[18:0], v3589[20:0]); // 3.0
    wire [13:0] v3590; shift_adder #(11, 14, 1, 1, 14, -1, 0) op_3590 (v1943[10:0], v1944[13:0], v3590[13:0]); // 3.0
    wire [24:0] v3591; shift_adder #(22, 19, 1, 1, 25, 6, 0) op_3591 (v1365[21:0], v1945[18:0], v3591[24:0]); // 3.0
    wire [13:0] v3592; shift_adder #(12, 13, 1, 1, 14, -2, 0) op_3592 (v1069[11:0], v1946[12:0], v3592[13:0]); // 3.0
    wire [26:0] v3593; shift_adder #(12, 15, 1, 1, 27, -15, 0) op_3593 (v1462[11:0], v1947[14:0], v3593[26:0]); // 3.0
    wire [12:0] v3594; shift_adder #(12, 13, 1, 1, 13, 0, 0) op_3594 (v1730[11:0], v1187[12:0], v3594[12:0]); // 3.0
    wire [11:0] v3595; shift_adder #(11, 11, 1, 1, 12, 0, 1) op_3595 (v1122[10:0], v400[10:0], v3595[11:0]); // 3.0
    wire [15:0] v3596; shift_adder #(12, 16, 1, 1, 16, -2, 0) op_3596 (v292[11:0], v1913[15:0], v3596[15:0]); // 3.0
    wire [24:0] v3597; shift_adder #(25, 12, 1, 1, 25, 11, 0) op_3597 (v1625[24:0], v873[11:0], v3597[24:0]); // 3.0
    wire [14:0] v3598; shift_adder #(14, 14, 1, 1, 15, 0, 0) op_3598 (v1250[13:0], v1522[13:0], v3598[14:0]); // 3.0
    wire [13:0] v3599; shift_adder #(12, 13, 1, 1, 14, -1, 0) op_3599 (v1948[11:0], v1949[12:0], v3599[13:0]); // 3.0
    wire [17:0] v3600; shift_adder #(16, 16, 1, 1, 18, 2, 0) op_3600 (v1525[15:0], v1950[15:0], v3600[17:0]); // 3.0
    wire [16:0] v3601; shift_adder #(11, 12, 1, 1, 17, 5, 1) op_3601 (v150[10:0], v1726[11:0], v3601[16:0]); // 3.0
    wire [15:0] v3602; shift_adder #(11, 13, 1, 1, 16, -5, 0) op_3602 (v518[10:0], v793[12:0], v3602[15:0]); // 3.0
    wire [14:0] v3603; shift_adder #(12, 12, 1, 1, 15, 3, 0) op_3603 (v854[11:0], v1951[11:0], v3603[14:0]); // 3.0
    wire [13:0] v3604; shift_adder #(12, 13, 1, 1, 14, 0, 0) op_3604 (v1865[11:0], v1097[12:0], v3604[13:0]); // 3.0
    wire [30:0] v3605; shift_adder #(12, 29, 1, 1, 31, -18, 0) op_3605 (v1025[11:0], v1952[28:0], v3605[30:0]); // 3.0
    wire [33:0] v3606; shift_adder #(13, 33, 1, 1, 34, -19, 0) op_3606 (v1263[12:0], v1953[32:0], v3606[33:0]); // 3.0
    wire [21:0] v3607; shift_adder #(17, 21, 1, 1, 22, -5, 0) op_3607 (v551[16:0], v1596[20:0], v3607[21:0]); // 3.0
    wire [22:0] v3608; shift_adder #(23, 11, 1, 1, 23, 11, 0) op_3608 (v1954[22:0], v961[10:0], v3608[22:0]); // 3.0
    wire [13:0] v3609; shift_adder #(13, 12, 1, 1, 14, 2, 0) op_3609 (v1955[12:0], v1956[11:0], v3609[13:0]); // 3.0
    wire [39:0] v3610; shift_adder #(13, 11, 1, 1, 40, 29, 1) op_3610 (v1021[12:0], v497[10:0], v3610[39:0]); // 3.0
    wire [12:0] v3611; shift_adder #(12, 12, 1, 1, 13, 1, 0) op_3611 (v1957[11:0], v1958[11:0], v3611[12:0]); // 3.0
    wire [14:0] v3612; shift_adder #(12, 12, 1, 1, 15, 2, 0) op_3612 (v924[11:0], v1649[11:0], v3612[14:0]); // 3.0
    wire [36:0] v3613; shift_adder #(36, 26, 1, 1, 37, 11, 0) op_3613 (v1959[35:0], v1449[25:0], v3613[36:0]); // 3.0
    wire [17:0] v3614; shift_adder #(11, 16, 1, 1, 18, -6, 0) op_3614 (v1960[10:0], v1961[15:0], v3614[17:0]); // 3.0
    wire [18:0] v3615; shift_adder #(12, 17, 1, 1, 19, -6, 0) op_3615 (v1511[11:0], v963[16:0], v3615[18:0]); // 3.0
    wire [14:0] v3616; shift_adder #(14, 12, 1, 1, 15, 1, 0) op_3616 (v1962[13:0], v1637[11:0], v3616[14:0]); // 3.0
    wire [13:0] v3617; shift_adder #(12, 12, 1, 1, 14, 1, 0) op_3617 (v1963[11:0], v1631[11:0], v3617[13:0]); // 3.0
    wire [15:0] v3618; shift_adder #(15, 11, 1, 1, 16, 3, 0) op_3618 (v1964[14:0], v1965[10:0], v3618[15:0]); // 3.0
    wire [18:0] v3619; shift_adder #(11, 19, 1, 1, 19, -2, 0) op_3619 (v259[10:0], v1966[18:0], v3619[18:0]); // 3.0
    wire [22:0] v3620; shift_adder #(21, 13, 1, 1, 23, 9, 0) op_3620 (v1144[20:0], v1967[12:0], v3620[22:0]); // 3.0
    wire [15:0] v3621; shift_adder #(8, 13, 1, 1, 16, 3, 0) op_3621 (v108[7:0], v883[12:0], v3621[15:0]); // 3.0
    wire [26:0] v3622; shift_adder #(26, 17, 1, 1, 27, 10, 0) op_3622 (v1882[25:0], v881[16:0], v3622[26:0]); // 3.0
    wire [24:0] v3623; shift_adder #(13, 23, 1, 1, 25, -11, 0) op_3623 (v1968[12:0], v1743[22:0], v3623[24:0]); // 3.0
    wire [22:0] v3624; shift_adder #(23, 13, 1, 1, 23, 5, 1) op_3624 (v1733[22:0], v1524[12:0], v3624[22:0]); // 3.0
    wire [17:0] v3625; shift_adder #(17, 15, 1, 1, 18, 3, 0) op_3625 (v1312[16:0], v1628[14:0], v3625[17:0]); // 3.0
    wire [25:0] v3626; shift_adder #(26, 25, 1, 1, 26, 0, 0) op_3626 (v988[25:0], v1935[24:0], v3626[25:0]); // 3.0
    wire [16:0] v3627; shift_adder #(16, 12, 1, 1, 17, 3, 0) op_3627 (v1969[15:0], v896[11:0], v3627[16:0]); // 3.0
    wire [17:0] v3628; shift_adder #(17, 13, 1, 1, 18, 3, 0) op_3628 (v1063[16:0], v818[12:0], v3628[17:0]); // 3.0
    wire [16:0] v3629; shift_adder #(13, 16, 1, 1, 17, -4, 0) op_3629 (v1970[12:0], v1414[15:0], v3629[16:0]); // 3.0
    wire [24:0] v3630; shift_adder #(23, 14, 1, 1, 25, 10, 0) op_3630 (v1971[22:0], v1972[13:0], v3630[24:0]); // 3.0
    wire [17:0] v3631; shift_adder #(12, 14, 1, 1, 18, -6, 0) op_3631 (v586[11:0], v1973[13:0], v3631[17:0]); // 3.0
    wire [23:0] v3632; shift_adder #(24, 13, 1, 1, 24, 10, 0) op_3632 (v1418[23:0], v1974[12:0], v3632[23:0]); // 3.0
    wire [20:0] v3633; shift_adder #(15, 21, 1, 1, 21, -4, 0) op_3633 (v1975[14:0], v1976[20:0], v3633[20:0]); // 3.0
    wire [20:0] v3634; shift_adder #(12, 19, 1, 1, 21, -8, 0) op_3634 (v1977[11:0], v1644[18:0], v3634[20:0]); // 3.0
    wire [17:0] v3635; shift_adder #(8, 18, 1, 1, 18, -6, 0) op_3635 (v99[7:0], v1978[17:0], v3635[17:0]); // 3.0
    wire [15:0] v3636; shift_adder #(14, 15, 1, 1, 16, -1, 0) op_3636 (v1979[13:0], v913[14:0], v3636[15:0]); // 3.0
    wire [17:0] v3637; shift_adder #(18, 12, 1, 1, 18, 4, 0) op_3637 (v789[17:0], v475[11:0], v3637[17:0]); // 3.0
    wire [21:0] v3638; shift_adder #(14, 21, 1, 1, 22, -6, 0) op_3638 (v1980[13:0], v1981[20:0], v3638[21:0]); // 3.0
    wire [19:0] v3639; shift_adder #(14, 20, 1, 1, 20, -5, 0) op_3639 (v1982[13:0], v1983[19:0], v3639[19:0]); // 3.0
    wire [19:0] v3640; shift_adder #(14, 20, 1, 1, 20, -3, 1) op_3640 (v1420[13:0], v1984[19:0], v3640[19:0]); // 3.0
    wire [14:0] v3641; shift_adder #(15, 11, 1, 1, 15, 0, 1) op_3641 (v1576[14:0], v821[10:0], v3641[14:0]); // 3.0
    wire [22:0] v3642; shift_adder #(19, 22, 1, 1, 23, -3, 0) op_3642 (v1565[18:0], v804[21:0], v3642[22:0]); // 3.0
    wire [12:0] v3643; shift_adder #(12, 12, 1, 1, 13, 0, 0) op_3643 (v1573[11:0], v1940[11:0], v3643[12:0]); // 3.0
    wire [29:0] v3644; shift_adder #(24, 28, 1, 1, 30, -6, 0) op_3644 (v1470[23:0], v1771[27:0], v3644[29:0]); // 3.0
    wire [18:0] v3645; shift_adder #(18, 13, 1, 1, 19, 5, 0) op_3645 (v1502[17:0], v1985[12:0], v3645[18:0]); // 3.0
    wire [13:0] v3646; shift_adder #(12, 13, 1, 1, 14, -1, 0) op_3646 (v1986[11:0], v1397[12:0], v3646[13:0]); // 3.0
    wire [17:0] v3647; shift_adder #(18, 15, 1, 1, 18, 2, 0) op_3647 (v1987[17:0], v1499[14:0], v3647[17:0]); // 3.0
    wire [27:0] v3648; shift_adder #(22, 27, 1, 1, 28, -5, 0) op_3648 (v1988[21:0], v1989[26:0], v3648[27:0]); // 3.0
    wire [33:0] v3649; shift_adder #(34, 12, 1, 1, 34, 21, 0) op_3649 (v1597[33:0], v1990[11:0], v3649[33:0]); // 3.0
    wire [12:0] v3650; shift_adder #(13, 11, 1, 1, 13, 0, 0) op_3650 (v1359[12:0], v772[10:0], v3650[12:0]); // 3.0
    wire [17:0] v3651; shift_adder #(17, 13, 1, 1, 18, 3, 0) op_3651 (v1991[16:0], v1992[12:0], v3651[17:0]); // 3.0
    wire [15:0] v3652; shift_adder #(13, 14, 1, 1, 16, -2, 0) op_3652 (v880[12:0], v1300[13:0], v3652[15:0]); // 3.0
    wire [23:0] v3653; shift_adder #(12, 23, 1, 1, 24, 1, 0) op_3653 (v1136[11:0], v1993[22:0], v3653[23:0]); // 3.0
    wire [13:0] v3654; shift_adder #(12, 13, 1, 1, 14, -2, 1) op_3654 (v452[11:0], v1404[12:0], v3654[13:0]); // 3.0
    wire [15:0] v3655; shift_adder #(13, 14, 1, 1, 16, -2, 0) op_3655 (v883[12:0], v1927[13:0], v3655[15:0]); // 3.0
    wire [30:0] v3656; shift_adder #(23, 29, 1, 1, 31, -8, 0) op_3656 (v1797[22:0], v1994[28:0], v3656[30:0]); // 3.0
    wire [16:0] v3657; shift_adder #(12, 16, 1, 1, 17, -4, 0) op_3657 (v1995[11:0], v1827[15:0], v3657[16:0]); // 3.0
    wire [32:0] v3658; shift_adder #(12, 10, 1, 1, 33, 23, 1) op_3658 (v1996[11:0], v516[9:0], v3658[32:0]); // 3.0
    wire [18:0] v3659; shift_adder #(13, 19, 1, 1, 19, -5, 0) op_3659 (v1677[12:0], v1900[18:0], v3659[18:0]); // 3.0
    wire [13:0] v3660; shift_adder #(13, 13, 1, 1, 14, -1, 0) op_3660 (v1997[12:0], v1998[12:0], v3660[13:0]); // 3.0
    wire [19:0] v3661; shift_adder #(12, 19, 1, 1, 20, -6, 0) op_3661 (v1199[11:0], v1999[18:0], v3661[19:0]); // 3.0
    wire [13:0] v3662; shift_adder #(13, 14, 1, 1, 14, 0, 0) op_3662 (v793[12:0], v1135[13:0], v3662[13:0]); // 3.0
    wire [13:0] v3663; shift_adder #(12, 13, 1, 1, 14, 0, 0) op_3663 (v1262[11:0], v915[12:0], v3663[13:0]); // 3.0
    wire [13:0] v3664; shift_adder #(12, 12, 1, 1, 14, -2, 0) op_3664 (v2000[11:0], v2001[11:0], v3664[13:0]); // 3.0
    wire [19:0] v3665; shift_adder #(16, 17, 1, 1, 20, -4, 0) op_3665 (v1020[15:0], v1146[16:0], v3665[19:0]); // 3.0
    wire [14:0] v3666; shift_adder #(11, 13, 1, 1, 15, -4, 1) op_3666 (v386[10:0], v1446[12:0], v3666[14:0]); // 3.0
    wire [15:0] v3667; shift_adder #(12, 13, 1, 1, 16, -4, 0) op_3667 (v1631[11:0], v2002[12:0], v3667[15:0]); // 3.0
    wire [15:0] v3668; shift_adder #(14, 13, 1, 1, 16, 2, 0) op_3668 (v1545[13:0], v1336[12:0], v3668[15:0]); // 3.0
    wire [14:0] v3669; shift_adder #(15, 12, 1, 1, 15, 2, 0) op_3669 (v2003[14:0], v2004[11:0], v3669[14:0]); // 3.0
    wire [24:0] v3670; shift_adder #(11, 25, 1, 1, 25, -6, 0) op_3670 (v140[10:0], v1875[24:0], v3670[24:0]); // 3.0
    wire [17:0] v3671; shift_adder #(12, 18, 1, 1, 18, 0, 1) op_3671 (v1398[11:0], v938[17:0], v3671[17:0]); // 3.0
    wire [24:0] v3672; shift_adder #(8, 15, 1, 1, 25, -16, 0) op_3672 (v109[7:0], v2005[14:0], v3672[24:0]); // 3.0
    wire [26:0] v3673; shift_adder #(27, 14, 1, 1, 27, 11, 0) op_3673 (v1579[26:0], v1516[13:0], v3673[26:0]); // 3.0
    wire [17:0] v3674; shift_adder #(17, 12, 1, 1, 18, 5, 0) op_3674 (v1526[16:0], v1443[11:0], v3674[17:0]); // 3.0
    wire [16:0] v3675; shift_adder #(13, 16, 1, 1, 17, -3, 0) op_3675 (v859[12:0], v1541[15:0], v3675[16:0]); // 3.0
    wire [22:0] v3676; shift_adder #(16, 23, 1, 1, 23, -5, 0) op_3676 (v1238[15:0], v811[22:0], v3676[22:0]); // 3.0
    wire [23:0] v3677; shift_adder #(24, 17, 1, 1, 24, 4, 0) op_3677 (v2006[23:0], v2007[16:0], v3677[23:0]); // 3.0
    wire [17:0] v3678; shift_adder #(18, 14, 1, 1, 18, 3, 0) op_3678 (v1692[17:0], v2008[13:0], v3678[17:0]); // 3.0
    wire [15:0] v3679; shift_adder #(13, 13, 1, 1, 16, 3, 0) op_3679 (v149[12:0], v1074[12:0], v3679[15:0]); // 3.0
    wire [24:0] v3680; shift_adder #(8, 25, 1, 1, 25, -9, 1) op_3680 (v123[7:0], v2009[24:0], v3680[24:0]); // 3.0
    wire [15:0] v3681; shift_adder #(13, 16, 1, 1, 16, -2, 0) op_3681 (v2010[12:0], v1717[15:0], v3681[15:0]); // 3.0
    wire [29:0] v3682; shift_adder #(29, 14, 1, 1, 30, 15, 0) op_3682 (v850[28:0], v2011[13:0], v3682[29:0]); // 3.0
    wire [29:0] v3683; shift_adder #(30, 11, 1, 1, 30, 17, 0) op_3683 (v1239[29:0], v1492[10:0], v3683[29:0]); // 3.0
    wire [30:0] v3684; shift_adder #(30, 17, 1, 1, 31, 13, 0) op_3684 (v2012[29:0], v1809[16:0], v3684[30:0]); // 3.0
    wire [13:0] v3685; shift_adder #(13, 12, 1, 1, 14, 2, 0) op_3685 (v1482[12:0], v1413[11:0], v3685[13:0]); // 3.0
    wire [20:0] v3686; shift_adder #(15, 21, 1, 1, 21, -5, 0) op_3686 (v1439[14:0], v1596[20:0], v3686[20:0]); // 3.0
    wire [15:0] v3687; shift_adder #(14, 15, 1, 1, 16, -2, 1) op_3687 (v555[13:0], v1401[14:0], v3687[15:0]); // 3.0
    wire [19:0] v3688; shift_adder #(18, 13, 1, 1, 20, 7, 0) op_3688 (v2013[17:0], v2014[12:0], v3688[19:0]); // 3.0
    wire [15:0] v3689; shift_adder #(11, 15, 1, 1, 16, -4, 0) op_3689 (v1358[10:0], v2015[14:0], v3689[15:0]); // 3.0
    wire [16:0] v3690; shift_adder #(16, 12, 1, 1, 17, 5, 0) op_3690 (v849[15:0], v1259[11:0], v3690[16:0]); // 3.0
    wire [14:0] v3691; shift_adder #(13, 15, 1, 1, 15, -1, 0) op_3691 (v1263[12:0], v2016[14:0], v3691[14:0]); // 3.0
    wire [18:0] v3692; shift_adder #(17, 15, 1, 1, 19, 3, 0) op_3692 (v1231[16:0], v1053[14:0], v3692[18:0]); // 3.0
    wire [12:0] v3693; shift_adder #(11, 12, 1, 1, 13, -1, 0) op_3693 (v885[10:0], v2017[11:0], v3693[12:0]); // 3.0
    wire [12:0] v3694; shift_adder #(12, 12, 1, 1, 13, 0, 0) op_3694 (v936[11:0], v2019[11:0], v3694[12:0]); // 3.0
    wire [16:0] v3695; shift_adder #(15, 12, 1, 1, 17, 4, 0) op_3695 (v2020[14:0], v1171[11:0], v3695[16:0]); // 3.0
    wire [14:0] v3696; shift_adder #(8, 13, 1, 1, 15, 2, 0) op_3696 (v111[7:0], v1034[12:0], v3696[14:0]); // 3.0
    wire [24:0] v3697; shift_adder #(24, 19, 1, 1, 25, 5, 0) op_3697 (v1734[23:0], v2021[18:0], v3697[24:0]); // 3.0
    wire [22:0] v3698; shift_adder #(12, 15, 1, 1, 23, 8, 1) op_3698 (v452[11:0], v2022[14:0], v3698[22:0]); // 3.0
    wire [18:0] v3699; shift_adder #(18, 18, 1, 1, 19, 0, 0) op_3699 (v1987[17:0], v1005[17:0], v3699[18:0]); // 3.0
    wire [21:0] v3700; shift_adder #(12, 22, 1, 1, 22, -5, 0) op_3700 (v1370[11:0], v2023[21:0], v3700[21:0]); // 3.0
    wire [12:0] v3701; shift_adder #(8, 13, 1, 1, 13, -1, 0) op_3701 (v107[7:0], v1030[12:0], v3701[12:0]); // 3.0
    wire [15:0] v3702; shift_adder #(13, 12, 1, 1, 16, 4, 0) op_3702 (v2024[12:0], v1234[11:0], v3702[15:0]); // 3.0
    wire [25:0] v3703; shift_adder #(18, 11, 1, 1, 26, -8, 0) op_3703 (v2025[17:0], v954[10:0], v3703[25:0]); // 3.0
    wire [26:0] v3704; shift_adder #(26, 15, 1, 1, 27, 11, 0) op_3704 (v979[25:0], v1038[14:0], v3704[26:0]); // 3.0
    wire [17:0] v3705; shift_adder #(16, 17, 1, 1, 18, -1, 0) op_3705 (v927[15:0], v952[16:0], v3705[17:0]); // 3.0
    wire [15:0] v3706; shift_adder #(11, 16, 1, 1, 16, -1, 1) op_3706 (v217[10:0], v1525[15:0], v3706[15:0]); // 3.0
    wire [25:0] v3707; shift_adder #(16, 25, 1, 1, 26, -9, 0) op_3707 (v1531[15:0], v2026[24:0], v3707[25:0]); // 3.0
    wire [22:0] v3708; shift_adder #(16, 12, 1, 1, 23, -7, 0) op_3708 (v426[15:0], v2027[11:0], v3708[22:0]); // 3.0
    wire [33:0] v3709; shift_adder #(33, 14, 1, 1, 34, 19, 0) op_3709 (v1441[32:0], v2028[13:0], v3709[33:0]); // 3.0
    wire [28:0] v3710; shift_adder #(28, 15, 1, 1, 29, 13, 0) op_3710 (v2029[27:0], v894[14:0], v3710[28:0]); // 3.0
    wire [13:0] v3711; shift_adder #(11, 13, 1, 1, 14, -2, 0) op_3711 (v153[10:0], v803[12:0], v3711[13:0]); // 3.0
    wire [23:0] v3712; shift_adder #(23, 12, 1, 1, 24, 11, 0) op_3712 (v1648[22:0], v2030[11:0], v3712[23:0]); // 3.0
    wire [16:0] v3713; shift_adder #(12, 13, 1, 1, 17, -5, 0) op_3713 (v1082[11:0], v2031[12:0], v3713[16:0]); // 3.0
    wire [23:0] v3714; shift_adder #(15, 22, 1, 1, 24, -9, 0) op_3714 (v1919[14:0], v2032[21:0], v3714[23:0]); // 3.0
    wire [26:0] v3715; shift_adder #(15, 19, 1, 1, 27, 8, 0) op_3715 (v905[14:0], v2034[18:0], v3715[26:0]); // 3.0
    wire [14:0] v3716; shift_adder #(12, 13, 1, 1, 15, 1, 0) op_3716 (v848[11:0], v2035[12:0], v3716[14:0]); // 3.0
    wire [15:0] v3717; shift_adder #(11, 13, 1, 1, 16, -4, 0) op_3717 (v1306[10:0], v1247[12:0], v3717[15:0]); // 3.0
    wire [17:0] v3718; shift_adder #(18, 14, 1, 1, 18, 3, 0) op_3718 (v1778[17:0], v2036[13:0], v3718[17:0]); // 3.0
    wire [17:0] v3719; shift_adder #(17, 11, 1, 1, 18, -1, 0) op_3719 (v143[16:0], v1943[10:0], v3719[17:0]); // 3.0
    wire [20:0] v3720; shift_adder #(12, 12, 1, 1, 21, 9, 1) op_3720 (v457[11:0], v1147[11:0], v3720[20:0]); // 3.0
    wire [15:0] v3721; shift_adder #(16, 15, 1, 1, 16, 0, 0) op_3721 (v1064[15:0], v2037[14:0], v3721[15:0]); // 3.0
    wire [21:0] v3722; shift_adder #(21, 12, 1, 1, 22, 9, 0) op_3722 (v2038[20:0], v2039[11:0], v3722[21:0]); // 3.0
    wire [34:0] v3723; shift_adder #(14, 24, 1, 1, 35, -21, 0) op_3723 (v2040[13:0], v2041[23:0], v3723[34:0]); // 3.0
    wire [16:0] v3724; shift_adder #(16, 16, 1, 1, 17, 0, 0) op_3724 (v814[15:0], v1389[15:0], v3724[16:0]); // 3.0
    wire [27:0] v3725; shift_adder #(12, 14, 1, 1, 28, -16, 1) op_3725 (v159[11:0], v1002[13:0], v3725[27:0]); // 3.0
    wire [23:0] v3726; shift_adder #(22, 19, 1, 1, 24, 4, 0) op_3726 (v2042[21:0], v1830[18:0], v3726[23:0]); // 3.0
    wire [13:0] v3727; shift_adder #(12, 11, 1, 1, 14, 2, 0) op_3727 (v1585[11:0], v1905[10:0], v3727[13:0]); // 3.0
    wire [14:0] v3728; shift_adder #(14, 14, 1, 1, 15, 0, 0) op_3728 (v1317[13:0], v1381[13:0], v3728[14:0]); // 3.0
    wire [16:0] v3729; shift_adder #(12, 15, 1, 1, 17, -4, 0) op_3729 (v2043[11:0], v2044[14:0], v3729[16:0]); // 3.0
    wire [24:0] v3730; shift_adder #(25, 14, 1, 1, 25, 10, 0) op_3730 (v1544[24:0], v2045[13:0], v3730[24:0]); // 3.0
    wire [20:0] v3731; shift_adder #(12, 15, 1, 1, 21, 6, 0) op_3731 (v1069[11:0], v904[14:0], v3731[20:0]); // 3.0
    wire [18:0] v3732; shift_adder #(15, 18, 1, 1, 19, -3, 0) op_3732 (v2046[14:0], v2047[17:0], v3732[18:0]); // 3.0
    wire [16:0] v3733; shift_adder #(8, 14, 1, 1, 17, -8, 0) op_3733 (v84[7:0], v2048[13:0], v3733[16:0]); // 3.0
    wire [19:0] v3734; shift_adder #(19, 14, 1, 1, 20, 4, 0) op_3734 (v1626[18:0], v2049[13:0], v3734[19:0]); // 3.0
    wire [36:0] v3735; shift_adder #(21, 36, 1, 1, 37, -16, 0) op_3735 (v1090[20:0], v2050[35:0], v3735[36:0]); // 3.0
    wire [30:0] v3736; shift_adder #(13, 30, 1, 1, 31, -17, 0) op_3736 (v1404[12:0], v1442[29:0], v3736[30:0]); // 3.0
    wire [22:0] v3737; shift_adder #(11, 15, 1, 1, 23, -12, 0) op_3737 (v297[10:0], v1205[14:0], v3737[22:0]); // 3.0
    wire [14:0] v3738; shift_adder #(11, 15, 1, 1, 15, -2, 0) op_3738 (v238[10:0], v1272[14:0], v3738[14:0]); // 3.0
    wire [23:0] v3739; shift_adder #(23, 12, 1, 1, 24, 11, 0) op_3739 (v980[22:0], v1259[11:0], v3739[23:0]); // 3.0
    wire [32:0] v3740; shift_adder #(11, 13, 1, 1, 33, 20, 1) op_3740 (v2051[10:0], v654[12:0], v3740[32:0]); // 3.0
    wire [29:0] v3741; shift_adder #(29, 19, 1, 1, 30, 10, 0) op_3741 (v1952[28:0], v2052[18:0], v3741[29:0]); // 3.0
    wire [15:0] v3742; shift_adder #(15, 11, 1, 1, 16, 3, 0) op_3742 (v2053[14:0], v2054[10:0], v3742[15:0]); // 3.0
    wire [19:0] v3743; shift_adder #(20, 14, 1, 1, 20, 5, 0) op_3743 (v2055[19:0], v2056[13:0], v3743[19:0]); // 3.0
    wire [37:0] v3744; shift_adder #(35, 37, 1, 1, 38, -1, 0) op_3744 (v2057[34:0], v2058[36:0], v3744[37:0]); // 3.0
    wire [13:0] v3745; shift_adder #(12, 12, 1, 1, 14, -2, 0) op_3745 (v1370[11:0], v2059[11:0], v3745[13:0]); // 3.0
    wire [15:0] v3746; shift_adder #(16, 13, 1, 1, 16, 1, 0) op_3746 (v1719[15:0], v833[12:0], v3746[15:0]); // 3.0
    wire [16:0] v3747; shift_adder #(13, 15, 1, 1, 17, -3, 0) op_3747 (v1041[12:0], v2060[14:0], v3747[16:0]); // 3.0
    wire [14:0] v3748; shift_adder #(12, 13, 1, 1, 15, -3, 0) op_3748 (v2061[11:0], v2062[12:0], v3748[14:0]); // 3.0
    wire [13:0] v3749; shift_adder #(12, 13, 1, 1, 14, -2, 0) op_3749 (v2063[11:0], v1078[12:0], v3749[13:0]); // 3.0
    wire [13:0] v3750; shift_adder #(12, 13, 1, 1, 14, 0, 0) op_3750 (v2064[11:0], v2065[12:0], v3750[13:0]); // 3.0
    wire [20:0] v3751; shift_adder #(11, 13, 1, 1, 21, 8, 1) op_3751 (v420[10:0], v1029[12:0], v3751[20:0]); // 3.0
    wire [17:0] v3752; shift_adder #(15, 16, 1, 1, 18, -3, 0) op_3752 (v1186[14:0], v1452[15:0], v3752[17:0]); // 3.0
    wire [18:0] v3753; shift_adder #(19, 13, 1, 1, 19, 3, 0) op_3753 (v1830[18:0], v1097[12:0], v3753[18:0]); // 3.0
    wire [17:0] v3754; shift_adder #(13, 17, 1, 1, 18, -4, 0) op_3754 (v2066[12:0], v1157[16:0], v3754[17:0]); // 3.0
    wire [19:0] v3755; shift_adder #(8, 12, 1, 1, 20, 8, 1) op_3755 (v73[7:0], v1555[11:0], v3755[19:0]); // 3.0
    wire [15:0] v3756; shift_adder #(14, 15, 1, 1, 16, 1, 0) op_3756 (v2067[13:0], v2068[14:0], v3756[15:0]); // 3.0
    wire [21:0] v3757; shift_adder #(11, 12, 1, 1, 22, 10, 1) op_3757 (v293[10:0], v1408[11:0], v3757[21:0]); // 3.0
    wire [20:0] v3758; shift_adder #(17, 18, 1, 1, 21, -4, 0) op_3758 (v2069[16:0], v1510[17:0], v3758[20:0]); // 3.0
    wire [21:0] v3759; shift_adder #(21, 15, 1, 1, 22, 6, 0) op_3759 (v2070[20:0], v1947[14:0], v3759[21:0]); // 3.0
    wire [16:0] v3760; shift_adder #(16, 15, 1, 1, 17, -1, 0) op_3760 (v1088[15:0], v1832[14:0], v3760[16:0]); // 3.0
    wire [22:0] v3761; shift_adder #(12, 19, 1, 1, 23, -11, 0) op_3761 (v202[11:0], v1830[18:0], v3761[22:0]); // 3.0
    wire [14:0] v3762; shift_adder #(12, 14, 1, 1, 15, -2, 0) op_3762 (v2071[11:0], v1834[13:0], v3762[14:0]); // 3.0
    wire [12:0] v3763; shift_adder #(12, 12, 1, 1, 13, 0, 0) op_3763 (v2072[11:0], v1612[11:0], v3763[12:0]); // 3.0
    wire [19:0] v3764; shift_adder #(15, 20, 1, 1, 20, -3, 0) op_3764 (v2073[14:0], v2074[19:0], v3764[19:0]); // 3.0
    wire [15:0] v3765; shift_adder #(8, 16, 1, 1, 16, -6, 0) op_3765 (v83[7:0], v1682[15:0], v3765[15:0]); // 3.0
    wire [23:0] v3766; shift_adder #(21, 24, 1, 1, 24, -1, 0) op_3766 (v1520[20:0], v780[23:0], v3766[23:0]); // 3.0
    wire [28:0] v3767; shift_adder #(28, 28, 1, 1, 29, 1, 0) op_3767 (v2029[27:0], v1504[27:0], v3767[28:0]); // 3.0
    wire [13:0] v3768; shift_adder #(9, 12, 1, 1, 14, -4, 1) op_3768 (v138[8:0], v1255[11:0], v3768[13:0]); // 3.0
    wire [26:0] v3769; shift_adder #(11, 13, 1, 1, 27, 14, 0) op_3769 (v237[10:0], v859[12:0], v3769[26:0]); // 3.0
    wire [24:0] v3770; shift_adder #(9, 14, 1, 1, 25, -15, 0) op_3770 (v395[8:0], v2075[13:0], v3770[24:0]); // 3.0
    wire [16:0] v3771; shift_adder #(13, 14, 1, 1, 17, -3, 0) op_3771 (v1599[12:0], v2076[13:0], v3771[16:0]); // 3.0
    wire [13:0] v3772; shift_adder #(12, 13, 1, 1, 14, 0, 0) op_3772 (v2077[11:0], v2078[12:0], v3772[13:0]); // 3.0
    wire [14:0] v3773; shift_adder #(15, 13, 1, 1, 15, 1, 0) op_3773 (v2079[14:0], v1782[12:0], v3773[14:0]); // 3.0
    wire [19:0] v3774; shift_adder #(19, 12, 1, 1, 20, 7, 0) op_3774 (v1217[18:0], v1570[11:0], v3774[19:0]); // 3.0
    wire [16:0] v3775; shift_adder #(16, 11, 1, 1, 17, 4, 0) op_3775 (v2080[15:0], v1711[10:0], v3775[16:0]); // 3.0
    wire [20:0] v3776; shift_adder #(19, 16, 1, 1, 21, 5, 0) op_3776 (v782[18:0], v959[15:0], v3776[20:0]); // 3.0
    wire [19:0] v3777; shift_adder #(16, 13, 1, 1, 20, -4, 0) op_3777 (v1620[15:0], v790[12:0], v3777[19:0]); // 3.0
    wire [14:0] v3778; shift_adder #(14, 13, 1, 1, 15, -1, 0) op_3778 (v1394[13:0], v2081[12:0], v3778[14:0]); // 3.0
    wire [20:0] v3779; shift_adder #(21, 14, 1, 1, 21, 4, 0) op_3779 (v907[20:0], v2082[13:0], v3779[20:0]); // 3.0
    wire [13:0] v3780; shift_adder #(12, 13, 1, 1, 14, 0, 0) op_3780 (v2083[11:0], v2084[12:0], v3780[13:0]); // 3.0
    wire [12:0] v3781; shift_adder #(12, 12, 1, 1, 13, 0, 0) op_3781 (v2085[11:0], v2086[11:0], v3781[12:0]); // 3.0
    wire [31:0] v3782; shift_adder #(18, 31, 1, 1, 32, -13, 0) op_3782 (v1592[17:0], v2087[30:0], v3782[31:0]); // 3.0
    wire [28:0] v3783; shift_adder #(8, 21, 1, 1, 29, 8, 0) op_3783 (v92[7:0], v1823[20:0], v3783[28:0]); // 3.0
    wire [22:0] v3784; shift_adder #(16, 22, 1, 1, 23, -7, 0) op_3784 (v2088[15:0], v2089[21:0], v3784[22:0]); // 3.0
    wire [19:0] v3785; shift_adder #(11, 13, 1, 1, 20, -9, 0) op_3785 (v341[10:0], v2090[12:0], v3785[19:0]); // 3.0
    wire [13:0] v3786; shift_adder #(13, 14, 1, 1, 14, 0, 0) op_3786 (v1230[12:0], v2091[13:0], v3786[13:0]); // 3.0
    wire [34:0] v3787; shift_adder #(12, 17, 1, 1, 35, 18, 1) op_3787 (v1555[11:0], v414[16:0], v3787[34:0]); // 3.0
    wire [34:0] v3788; shift_adder #(17, 35, 1, 1, 35, -7, 1) op_3788 (v1291[16:0], v2092[34:0], v3788[34:0]); // 3.0
    wire [20:0] v3789; shift_adder #(12, 12, 1, 1, 21, 9, 1) op_3789 (v408[11:0], v2072[11:0], v3789[20:0]); // 3.0
    wire [14:0] v3790; shift_adder #(13, 13, 1, 1, 15, 2, 0) op_3790 (v898[12:0], v1328[12:0], v3790[14:0]); // 3.0
    wire [35:0] v3791; shift_adder #(17, 12, 1, 1, 36, -19, 1) op_3791 (v2093[16:0], v2094[11:0], v3791[35:0]); // 3.0
    wire [15:0] v3792; shift_adder #(11, 15, 1, 1, 16, -4, 0) op_3792 (v2095[10:0], v2060[14:0], v3792[15:0]); // 3.0
    wire [28:0] v3793; shift_adder #(24, 28, 1, 1, 29, -4, 0) op_3793 (v2096[23:0], v2097[27:0], v3793[28:0]); // 3.0
    wire [16:0] v3794; shift_adder #(12, 17, 1, 1, 17, -4, 0) op_3794 (v447[11:0], v1700[16:0], v3794[16:0]); // 3.0
    wire [22:0] v3795; shift_adder #(14, 13, 1, 1, 23, -9, 1) op_3795 (v1162[13:0], v2098[12:0], v3795[22:0]); // 3.0
    wire [15:0] v3796; shift_adder #(15, 13, 1, 1, 16, 2, 0) op_3796 (v2099[14:0], v2100[12:0], v3796[15:0]); // 3.0
    wire [15:0] v3797; shift_adder #(13, 14, 1, 1, 16, -3, 0) op_3797 (v817[12:0], v2101[13:0], v3797[15:0]); // 3.0
    wire [19:0] v3798; shift_adder #(8, 17, 1, 1, 20, 3, 0) op_3798 (v99[7:0], v783[16:0], v3798[19:0]); // 3.0
    wire [15:0] v3799; shift_adder #(12, 15, 1, 1, 16, -3, 0) op_3799 (v1529[11:0], v1473[14:0], v3799[15:0]); // 3.0
    wire [15:0] v3800; shift_adder #(15, 11, 1, 1, 16, 4, 0) op_3800 (v1904[14:0], v2102[10:0], v3800[15:0]); // 3.0
    wire [25:0] v3801; shift_adder #(26, 14, 1, 1, 26, 9, 0) op_3801 (v2103[25:0], v1973[13:0], v3801[25:0]); // 3.0
    wire [19:0] v3802; shift_adder #(11, 15, 1, 1, 20, -9, 1) op_3802 (v328[10:0], v1417[14:0], v3802[19:0]); // 3.0
    wire [12:0] v3803; shift_adder #(10, 12, 1, 1, 13, -2, 0) op_3803 (v2104[9:0], v973[11:0], v3803[12:0]); // 3.0
    wire [26:0] v3804; shift_adder #(19, 27, 1, 1, 27, -3, 1) op_3804 (v782[18:0], v1878[26:0], v3804[26:0]); // 3.0
    wire [24:0] v3805; shift_adder #(24, 15, 1, 1, 25, 9, 0) op_3805 (v1807[23:0], v1867[14:0], v3805[24:0]); // 3.0
    wire [27:0] v3806; shift_adder #(9, 15, 1, 1, 28, 13, 0) op_3806 (v403[8:0], v2105[14:0], v3806[27:0]); // 3.0
    wire [23:0] v3807; shift_adder #(14, 10, 1, 1, 24, -10, 1) op_3807 (v1250[13:0], v489[9:0], v3807[23:0]); // 3.0
    wire [21:0] v3808; shift_adder #(12, 13, 1, 1, 22, 9, 0) op_3808 (v151[11:0], v1346[12:0], v3808[21:0]); // 3.0
    wire [15:0] v3809; shift_adder #(16, 15, 1, 1, 16, 0, 0) op_3809 (v1717[15:0], v2106[14:0], v3809[15:0]); // 3.0
    wire [15:0] v3810; shift_adder #(15, 12, 1, 1, 16, 2, 0) op_3810 (v1828[14:0], v2107[11:0], v3810[15:0]); // 3.0
    wire [22:0] v3811; shift_adder #(14, 12, 1, 1, 23, 11, 0) op_3811 (v342[13:0], v2108[11:0], v3811[22:0]); // 3.0
    wire [23:0] v3812; shift_adder #(23, 15, 1, 1, 24, 8, 0) op_3812 (v1648[22:0], v2109[14:0], v3812[23:0]); // 3.0
    wire [21:0] v3813; shift_adder #(21, 13, 1, 1, 22, 9, 0) op_3813 (v777[20:0], v1227[12:0], v3813[21:0]); // 3.0
    wire [15:0] v3814; shift_adder #(13, 16, 1, 1, 16, -2, 0) op_3814 (v2010[12:0], v1620[15:0], v3814[15:0]); // 3.0
    wire [22:0] v3815; shift_adder #(15, 23, 1, 1, 23, -5, 0) op_3815 (v1285[14:0], v1323[22:0], v3815[22:0]); // 3.0
    wire [15:0] v3816; shift_adder #(14, 15, 1, 1, 16, 1, 0) op_3816 (v2110[13:0], v2111[14:0], v3816[15:0]); // 3.0
    wire [17:0] v3817; shift_adder #(17, 17, 1, 1, 18, -1, 0) op_3817 (v1700[16:0], v2112[16:0], v3817[17:0]); // 3.0
    wire [16:0] v3818; shift_adder #(12, 15, 1, 1, 17, -4, 0) op_3818 (v1694[11:0], v1833[14:0], v3818[16:0]); // 3.0
    wire [21:0] v3819; shift_adder #(16, 14, 1, 1, 22, 8, 0) op_3819 (v1525[15:0], v342[13:0], v3819[21:0]); // 3.0
    wire [15:0] v3820; shift_adder #(15, 14, 1, 1, 16, -1, 0) op_3820 (v2113[14:0], v2056[13:0], v3820[15:0]); // 3.0
    wire [23:0] v3821; shift_adder #(11, 23, 1, 1, 24, -12, 1) op_3821 (v211[10:0], v2114[22:0], v3821[23:0]); // 3.0
    wire [21:0] v3822; shift_adder #(20, 14, 1, 1, 22, 8, 0) op_3822 (v1334[19:0], v2115[13:0], v3822[21:0]); // 3.0
    wire [18:0] v3823; shift_adder #(15, 18, 1, 1, 19, 1, 1) op_3823 (v2117[14:0], v1032[17:0], v3823[18:0]); // 3.0
    wire [23:0] v3824; shift_adder #(20, 14, 1, 1, 24, -4, 0) op_3824 (v1652[19:0], v2118[13:0], v3824[23:0]); // 3.0
    wire [18:0] v3825; shift_adder #(11, 18, 1, 1, 19, -7, 0) op_3825 (v821[10:0], v2013[17:0], v3825[18:0]); // 3.0
    wire [19:0] v3826; shift_adder #(20, 14, 1, 1, 20, 5, 0) op_3826 (v841[19:0], v1749[13:0], v3826[19:0]); // 3.0
    wire [22:0] v3827; shift_adder #(22, 11, 1, 1, 23, 11, 0) op_3827 (v909[21:0], v772[10:0], v3827[22:0]); // 3.0
    wire [18:0] v3828; shift_adder #(19, 16, 1, 1, 19, 2, 0) op_3828 (v2119[18:0], v959[15:0], v3828[18:0]); // 3.0
    wire [21:0] v3829; shift_adder #(21, 12, 1, 1, 22, 9, 0) op_3829 (v2120[20:0], v1171[11:0], v3829[21:0]); // 3.0
    wire [29:0] v3830; shift_adder #(30, 12, 1, 1, 30, 15, 0) op_3830 (v2121[29:0], v1155[11:0], v3830[29:0]); // 3.0
    wire [15:0] v3831; shift_adder #(14, 11, 1, 1, 16, 5, 0) op_3831 (v2122[13:0], v2123[10:0], v3831[15:0]); // 3.0
    wire [36:0] v3832; shift_adder #(12, 35, 1, 1, 37, -24, 0) op_3832 (v2124[11:0], v2125[34:0], v3832[36:0]); // 3.0
    wire [14:0] v3833; shift_adder #(13, 14, 1, 1, 15, -1, 0) op_3833 (v2126[12:0], v1045[13:0], v3833[14:0]); // 3.0
    wire [13:0] v3834; shift_adder #(12, 12, 1, 1, 14, -1, 0) op_3834 (v1080[11:0], v1160[11:0], v3834[13:0]); // 3.0
    wire [14:0] v3835; shift_adder #(13, 14, 1, 1, 15, 1, 0) op_3835 (v2127[12:0], v1695[13:0], v3835[14:0]); // 3.0
    wire [32:0] v3836; shift_adder #(33, 19, 1, 1, 33, 13, 0) op_3836 (v2128[32:0], v1217[18:0], v3836[32:0]); // 3.0
    wire [37:0] v3837; shift_adder #(17, 13, 1, 1, 38, -21, 1) op_3837 (v1619[16:0], v877[12:0], v3837[37:0]); // 3.0
    wire [15:0] v3838; shift_adder #(11, 15, 1, 1, 16, -3, 0) op_3838 (v2129[10:0], v866[14:0], v3838[15:0]); // 3.0
    wire [14:0] v3839; shift_adder #(15, 12, 1, 1, 15, 1, 0) op_3839 (v913[14:0], v2130[11:0], v3839[14:0]); // 3.0
    wire [20:0] v3840; shift_adder #(15, 20, 1, 1, 21, -6, 0) op_3840 (v1536[14:0], v2131[19:0], v3840[20:0]); // 3.0
    wire [16:0] v3841; shift_adder #(13, 17, 1, 1, 17, -3, 0) op_3841 (v884[12:0], v1291[16:0], v3841[16:0]); // 3.0
    wire [20:0] v3842; shift_adder #(21, 14, 1, 1, 21, 5, 0) op_3842 (v1722[20:0], v1317[13:0], v3842[20:0]); // 3.0
    wire [14:0] v3843; shift_adder #(12, 13, 1, 1, 15, -2, 0) op_3843 (v1277[11:0], v2132[12:0], v3843[14:0]); // 3.0
    wire [14:0] v3844; shift_adder #(13, 14, 1, 1, 15, -2, 0) op_3844 (v2133[12:0], v2134[13:0], v3844[14:0]); // 3.0
    wire [14:0] v3845; shift_adder #(12, 13, 1, 1, 15, -2, 0) op_3845 (v1309[11:0], v1569[12:0], v3845[14:0]); // 3.0
    wire [14:0] v3846; shift_adder #(11, 14, 1, 1, 15, -3, 0) op_3846 (v1137[10:0], v1818[13:0], v3846[14:0]); // 3.0
    wire [15:0] v3847; shift_adder #(12, 12, 1, 1, 16, 3, 0) op_3847 (v1153[11:0], v2135[11:0], v3847[15:0]); // 3.0
    wire [14:0] v3848; shift_adder #(14, 12, 1, 1, 15, 1, 0) op_3848 (v2136[13:0], v2137[11:0], v3848[14:0]); // 3.0
    wire [17:0] v3849; shift_adder #(14, 11, 1, 1, 18, 7, 0) op_3849 (v1222[13:0], v1306[10:0], v3849[17:0]); // 3.0
    wire [25:0] v3850; shift_adder #(13, 26, 1, 1, 26, -12, 0) op_3850 (v1787[12:0], v2138[25:0], v3850[25:0]); // 3.0
    wire [22:0] v3851; shift_adder #(16, 22, 1, 1, 23, -6, 0) op_3851 (v1114[15:0], v1061[21:0], v3851[22:0]); // 3.0
    wire [15:0] v3852; shift_adder #(15, 12, 1, 1, 16, 3, 0) op_3852 (v779[14:0], v1259[11:0], v3852[15:0]); // 3.0
    wire [13:0] v3853; shift_adder #(10, 13, 1, 1, 14, -2, 1) op_3853 (v643[9:0], v1665[12:0], v3853[13:0]); // 3.0
    wire [18:0] v3854; shift_adder #(19, 13, 1, 1, 19, 5, 0) op_3854 (v1565[18:0], v2139[12:0], v3854[18:0]); // 3.0
    wire [25:0] v3855; shift_adder #(13, 26, 1, 1, 26, -12, 1) op_3855 (v985[12:0], v802[25:0], v3855[25:0]); // 3.0
    wire [18:0] v3856; shift_adder #(11, 18, 1, 1, 19, -6, 0) op_3856 (v772[10:0], v2140[17:0], v3856[18:0]); // 3.0
    wire [14:0] v3857; shift_adder #(11, 13, 1, 1, 15, 2, 1) op_3857 (v1284[10:0], v1696[12:0], v3857[14:0]); // 3.0
    wire [13:0] v3858; shift_adder #(12, 13, 1, 1, 14, -1, 0) op_3858 (v2043[11:0], v2141[12:0], v3858[13:0]); // 3.0
    wire [31:0] v3859; shift_adder #(32, 18, 1, 1, 32, 11, 0) op_3859 (v1896[31:0], v2142[17:0], v3859[31:0]); // 3.0
    wire [15:0] v3860; shift_adder #(14, 15, 1, 1, 16, -1, 0) op_3860 (v2143[13:0], v1254[14:0], v3860[15:0]); // 3.0
    wire [22:0] v3861; shift_adder #(22, 21, 1, 1, 23, 1, 0) op_3861 (v2144[21:0], v1714[20:0], v3861[22:0]); // 3.0
    wire [32:0] v3862; shift_adder #(33, 22, 1, 1, 33, 9, 0) op_3862 (v1876[32:0], v1855[21:0], v3862[32:0]); // 3.0
    wire [27:0] v3863; shift_adder #(18, 27, 1, 1, 28, -10, 0) op_3863 (v2145[17:0], v1476[26:0], v3863[27:0]); // 3.0
    wire [14:0] v3864; shift_adder #(14, 12, 1, 1, 15, 2, 0) op_3864 (v2146[13:0], v1309[11:0], v3864[14:0]); // 3.0
    wire [15:0] v3865; shift_adder #(13, 14, 1, 1, 16, 2, 0) op_3865 (v859[12:0], v1813[13:0], v3865[15:0]); // 3.0
    wire [25:0] v3866; shift_adder #(16, 16, 1, 1, 26, -10, 1) op_3866 (v426[15:0], v1447[15:0], v3866[25:0]); // 3.0
    wire [16:0] v3867; shift_adder #(15, 12, 1, 1, 17, 4, 0) op_3867 (v1577[14:0], v1511[11:0], v3867[16:0]); // 3.0
    wire [25:0] v3868; shift_adder #(15, 25, 1, 1, 26, -10, 0) op_3868 (v1066[14:0], v2009[24:0], v3868[25:0]); // 3.0
    wire [15:0] v3869; shift_adder #(15, 14, 1, 1, 16, 1, 0) op_3869 (v1351[14:0], v2147[13:0], v3869[15:0]); // 3.0
    wire [29:0] v3870; shift_adder #(8, 30, 1, 1, 30, -6, 0) op_3870 (v117[7:0], v2148[29:0], v3870[29:0]); // 3.0
    wire [14:0] v3871; shift_adder #(14, 15, 1, 1, 15, 0, 0) op_3871 (v1420[13:0], v993[14:0], v3871[14:0]); // 3.0
    wire [16:0] v3872; shift_adder #(11, 15, 1, 1, 17, 2, 1) op_3872 (v171[10:0], v2005[14:0], v3872[16:0]); // 3.0
    wire [20:0] v3873; shift_adder #(12, 21, 1, 1, 21, -1, 0) op_3873 (v292[11:0], v1714[20:0], v3873[20:0]); // 3.0
    wire [21:0] v3874; shift_adder #(21, 12, 1, 1, 22, 9, 0) op_3874 (v2149[20:0], v1277[11:0], v3874[21:0]); // 3.0
    wire [16:0] v3875; shift_adder #(16, 13, 1, 1, 17, 4, 0) op_3875 (v2150[15:0], v1783[12:0], v3875[16:0]); // 3.0
    wire [20:0] v3876; shift_adder #(8, 16, 1, 1, 21, 5, 1) op_3876 (v75[7:0], v1913[15:0], v3876[20:0]); // 3.0
    wire [26:0] v3877; shift_adder #(21, 27, 1, 1, 27, -3, 0) op_3877 (v2038[20:0], v930[26:0], v3877[26:0]); // 3.0
    wire [24:0] v3878; shift_adder #(24, 12, 1, 1, 25, 12, 0) op_3878 (v2151[23:0], v2152[11:0], v3878[24:0]); // 3.0
    wire [18:0] v3879; shift_adder #(19, 12, 1, 1, 19, 4, 1) op_3879 (v1195[18:0], v267[11:0], v3879[18:0]); // 3.0
    wire [28:0] v3880; shift_adder #(12, 29, 1, 1, 29, -15, 0) op_3880 (v1347[11:0], v2153[28:0], v3880[28:0]); // 3.0
    wire [34:0] v3881; shift_adder #(15, 12, 1, 1, 35, 23, 1) op_3881 (v1127[14:0], v629[11:0], v3881[34:0]); // 3.0
    wire [13:0] v3882; shift_adder #(12, 12, 1, 1, 14, -2, 0) op_3882 (v2154[11:0], v2039[11:0], v3882[13:0]); // 3.0
    wire [16:0] v3883; shift_adder #(17, 12, 1, 1, 17, 3, 0) op_3883 (v2155[16:0], v1436[11:0], v3883[16:0]); // 3.0
    wire [15:0] v3884; shift_adder #(12, 15, 1, 1, 16, -2, 0) op_3884 (v1689[11:0], v815[14:0], v3884[15:0]); // 3.0
    wire [16:0] v3885; shift_adder #(13, 17, 1, 1, 17, -2, 0) op_3885 (v2156[12:0], v2157[16:0], v3885[16:0]); // 3.0
    wire [16:0] v3886; shift_adder #(14, 16, 1, 1, 17, -2, 0) op_3886 (v1132[13:0], v1762[15:0], v3886[16:0]); // 3.0
    wire [15:0] v3887; shift_adder #(12, 15, 1, 1, 16, -2, 0) op_3887 (v2158[11:0], v2159[14:0], v3887[15:0]); // 3.0
    wire [12:0] v3888; shift_adder #(8, 12, 1, 1, 13, -3, 1) op_3888 (v90[7:0], v2033[11:0], v3888[12:0]); // 3.0
    wire [16:0] v3889; shift_adder #(16, 12, 1, 1, 17, 4, 0) op_3889 (v1472[15:0], v1379[11:0], v3889[16:0]); // 3.0
    wire [30:0] v3890; shift_adder #(16, 30, 1, 1, 31, -13, 0) op_3890 (v2160[15:0], v1369[29:0], v3890[30:0]); // 3.0
    wire [18:0] v3891; shift_adder #(15, 19, 1, 1, 19, -3, 0) op_3891 (v1006[14:0], v2161[18:0], v3891[18:0]); // 3.0
    wire [26:0] v3892; shift_adder #(27, 15, 1, 1, 27, 11, 0) op_3892 (v912[26:0], v1027[14:0], v3892[26:0]); // 3.0
    wire [23:0] v3893; shift_adder #(21, 24, 1, 1, 24, -2, 0) op_3893 (v943[20:0], v1487[23:0], v3893[23:0]); // 3.0
    wire [19:0] v3894; shift_adder #(19, 15, 1, 1, 20, 5, 0) op_3894 (v1966[18:0], v1964[14:0], v3894[19:0]); // 3.0
    wire [16:0] v3895; shift_adder #(15, 12, 1, 1, 17, 4, 0) op_3895 (v781[14:0], v2162[11:0], v3895[16:0]); // 3.0
    wire [34:0] v3896; shift_adder #(34, 18, 1, 1, 35, 17, 0) op_3896 (v2163[33:0], v770[17:0], v3896[34:0]); // 3.0
    wire [14:0] v3897; shift_adder #(11, 11, 1, 1, 15, -3, 0) op_3897 (v2164[10:0], v772[10:0], v3897[14:0]); // 3.0
    wire [34:0] v3898; shift_adder #(12, 35, 1, 1, 35, -22, 0) op_3898 (v2165[11:0], v2166[34:0], v3898[34:0]); // 3.0
    wire [13:0] v3899; shift_adder #(13, 12, 1, 1, 14, 1, 0) op_3899 (v2167[12:0], v2168[11:0], v3899[13:0]); // 3.0
    wire [18:0] v3900; shift_adder #(19, 17, 1, 1, 19, 0, 0) op_3900 (v1218[18:0], v2169[16:0], v3900[18:0]); // 3.0
    wire [16:0] v3901; shift_adder #(13, 16, 1, 1, 17, -4, 0) op_3901 (v1422[12:0], v1552[15:0], v3901[16:0]); // 3.0
    wire [14:0] v3902; shift_adder #(11, 14, 1, 1, 15, -3, 1) op_3902 (v353[10:0], v1162[13:0], v3902[14:0]); // 3.0
    wire [13:0] v3903; shift_adder #(12, 13, 1, 1, 14, -1, 0) op_3903 (v1604[11:0], v2170[12:0], v3903[13:0]); // 3.0
    wire [17:0] v3904; shift_adder #(11, 13, 1, 1, 18, 5, 0) op_3904 (v301[10:0], v2171[12:0], v3904[17:0]); // 3.0
    wire [19:0] v3905; shift_adder #(20, 18, 1, 1, 20, 1, 0) op_3905 (v2172[19:0], v1130[17:0], v3905[19:0]); // 3.0
    wire [12:0] v3906; shift_adder #(13, 12, 1, 1, 13, 0, 0) op_3906 (v915[12:0], v1031[11:0], v3906[12:0]); // 3.0
    wire [33:0] v3907; shift_adder #(33, 17, 1, 1, 34, 16, 0) op_3907 (v1060[32:0], v1804[16:0], v3907[33:0]); // 3.0
    wire [22:0] v3908; shift_adder #(11, 13, 1, 1, 23, -12, 1) op_3908 (v276[10:0], v1704[12:0], v3908[22:0]); // 3.0
    wire [20:0] v3909; shift_adder #(11, 20, 1, 1, 21, -9, 0) op_3909 (v954[10:0], v1844[19:0], v3909[20:0]); // 3.0
    wire [30:0] v3910; shift_adder #(29, 17, 1, 1, 31, 14, 0) op_3910 (v1653[28:0], v2173[16:0], v3910[30:0]); // 3.0
    wire [18:0] v3911; shift_adder #(19, 18, 1, 1, 19, 0, 0) op_3911 (v2034[18:0], v1235[17:0], v3911[18:0]); // 3.0
    wire [25:0] v3912; shift_adder #(20, 24, 1, 1, 26, -6, 0) op_3912 (v1302[19:0], v1839[23:0], v3912[25:0]); // 3.0
    wire [16:0] v3913; shift_adder #(13, 15, 1, 1, 17, -3, 0) op_3913 (v2174[12:0], v1473[14:0], v3913[16:0]); // 3.0
    wire [14:0] v3914; shift_adder #(12, 13, 1, 1, 15, -3, 0) op_3914 (v1103[11:0], v1422[12:0], v3914[14:0]); // 3.0
    wire [15:0] v3915; shift_adder #(12, 12, 1, 1, 16, 4, 0) op_3915 (v227[11:0], v1659[11:0], v3915[15:0]); // 3.0
    wire [22:0] v3916; shift_adder #(13, 21, 1, 1, 23, 2, 1) op_3916 (v654[12:0], v1976[20:0], v3916[22:0]); // 3.0
    wire [18:0] v3917; shift_adder #(11, 18, 1, 1, 19, -7, 0) op_3917 (v1636[10:0], v968[17:0], v3917[18:0]); // 3.0
    wire [15:0] v3918; shift_adder #(15, 12, 1, 1, 16, 2, 0) op_3918 (v2175[14:0], v1754[11:0], v3918[15:0]); // 3.0
    wire [15:0] v3919; shift_adder #(16, 13, 1, 1, 16, 1, 0) op_3919 (v1620[15:0], v1397[12:0], v3919[15:0]); // 3.0
    wire [15:0] v3920; shift_adder #(15, 15, 1, 1, 16, 0, 0) op_3920 (v840[14:0], v1738[14:0], v3920[15:0]); // 3.0
    wire [13:0] v3921; shift_adder #(13, 13, 1, 1, 14, 0, 0) op_3921 (v2176[12:0], v2177[12:0], v3921[13:0]); // 3.0
    wire [16:0] v3922; shift_adder #(17, 15, 1, 1, 17, 0, 0) op_3922 (v889[16:0], v1874[14:0], v3922[16:0]); // 3.0
    wire [13:0] v3923; shift_adder #(13, 11, 1, 1, 14, 2, 1) op_3923 (v1189[12:0], v1284[10:0], v3923[13:0]); // 3.0
    wire [19:0] v3924; shift_adder #(12, 13, 1, 1, 20, -8, 0) op_3924 (v174[11:0], v813[12:0], v3924[19:0]); // 3.0
    wire [14:0] v3925; shift_adder #(14, 13, 1, 1, 15, 1, 0) op_3925 (v2178[13:0], v859[12:0], v3925[14:0]); // 3.0
    wire [14:0] v3926; shift_adder #(12, 12, 1, 1, 15, 2, 0) op_3926 (v1436[11:0], v2179[11:0], v3926[14:0]); // 3.0
    wire [14:0] v3927; shift_adder #(12, 14, 1, 1, 15, -2, 0) op_3927 (v2180[11:0], v2040[13:0], v3927[14:0]); // 3.0
    wire [17:0] v3928; shift_adder #(11, 15, 1, 1, 18, 3, 0) op_3928 (v415[10:0], v1535[14:0], v3928[17:0]); // 3.0
    wire [23:0] v3929; shift_adder #(11, 24, 1, 1, 24, -12, 0) op_3929 (v1581[10:0], v2181[23:0], v3929[23:0]); // 3.0
    wire [28:0] v3930; shift_adder #(18, 29, 1, 1, 29, -8, 0) op_3930 (v2182[17:0], v812[28:0], v3930[28:0]); // 3.0
    wire [20:0] v3931; shift_adder #(10, 21, 1, 1, 21, -9, 0) op_3931 (v2183[9:0], v1216[20:0], v3931[20:0]); // 3.0
    wire [21:0] v3932; shift_adder #(13, 21, 1, 1, 22, -8, 0) op_3932 (v2184[12:0], v1191[20:0], v3932[21:0]); // 3.0
    wire [15:0] v3933; shift_adder #(16, 14, 1, 1, 16, 1, 0) op_3933 (v2185[15:0], v1813[13:0], v3933[15:0]); // 3.0
    wire [15:0] v3934; shift_adder #(14, 15, 1, 1, 16, -1, 0) op_3934 (v2186[13:0], v1861[14:0], v3934[15:0]); // 3.0
    wire [17:0] v3935; shift_adder #(17, 11, 1, 1, 18, 6, 0) op_3935 (v2187[16:0], v1161[10:0], v3935[17:0]); // 3.0
    wire [25:0] v3936; shift_adder #(26, 12, 1, 1, 26, 12, 0) op_3936 (v1791[25:0], v2188[11:0], v3936[25:0]); // 3.0
    wire [15:0] v3937; shift_adder #(12, 15, 1, 1, 16, -4, 0) op_3937 (v1372[11:0], v922[14:0], v3937[15:0]); // 3.0
    wire [30:0] v3938; shift_adder #(14, 9, 1, 1, 31, 21, 1) op_3938 (v842[13:0], v663[8:0], v3938[30:0]); // 3.0
    wire [14:0] v3939; shift_adder #(8, 15, 1, 1, 15, 0, 1) op_3939 (v120[7:0], v1038[14:0], v3939[14:0]); // 3.0
    wire [16:0] v3940; shift_adder #(13, 15, 1, 1, 17, -4, 0) op_3940 (v892[12:0], v2189[14:0], v3940[16:0]); // 3.0
    wire [13:0] v3941; shift_adder #(12, 13, 1, 1, 14, 0, 0) op_3941 (v2190[11:0], v996[12:0], v3941[13:0]); // 3.0
    wire [15:0] v3942; shift_adder #(12, 14, 1, 1, 16, -3, 0) op_3942 (v1188[11:0], v1623[13:0], v3942[15:0]); // 3.0
    wire [34:0] v3943; shift_adder #(12, 33, 1, 1, 35, -23, 0) op_3943 (v820[11:0], v1051[32:0], v3943[34:0]); // 3.0
    wire [37:0] v3944; shift_adder #(36, 21, 1, 1, 38, 17, 0) op_3944 (v2191[35:0], v1040[20:0], v3944[37:0]); // 3.0
    wire [17:0] v3945; shift_adder #(13, 17, 1, 1, 18, -4, 0) op_3945 (v1021[12:0], v895[16:0], v3945[17:0]); // 3.0
    wire [15:0] v3946; shift_adder #(15, 13, 1, 1, 16, 2, 0) op_3946 (v2189[14:0], v2192[12:0], v3946[15:0]); // 3.0
    wire [35:0] v3947; shift_adder #(19, 11, 1, 1, 36, -17, 1) op_3947 (v2193[18:0], v2194[10:0], v3947[35:0]); // 3.0
    wire [13:0] v3948; shift_adder #(12, 11, 1, 1, 14, -1, 0) op_3948 (v1276[11:0], v2195[10:0], v3948[13:0]); // 3.0
    wire [18:0] v3949; shift_adder #(18, 19, 1, 1, 19, 0, 1) op_3949 (v2013[17:0], v1945[18:0], v3949[18:0]); // 3.0
    wire [23:0] v3950; shift_adder #(24, 16, 1, 1, 24, 7, 0) op_3950 (v2151[23:0], v1913[15:0], v3950[23:0]); // 3.0
    wire [13:0] v3951; shift_adder #(12, 12, 1, 1, 14, -1, 0) op_3951 (v2027[11:0], v1276[11:0], v3951[13:0]); // 3.0
    wire [19:0] v3952; shift_adder #(16, 20, 1, 1, 20, -1, 0) op_3952 (v1114[15:0], v1400[19:0], v3952[19:0]); // 3.0
    wire [18:0] v3953; shift_adder #(13, 17, 1, 1, 19, -5, 0) op_3953 (v2196[12:0], v890[16:0], v3953[18:0]); // 3.0
    wire [19:0] v3954; shift_adder #(19, 17, 1, 1, 20, 3, 0) op_3954 (v2197[18:0], v2198[16:0], v3954[19:0]); // 3.0
    wire [14:0] v3955; shift_adder #(11, 14, 1, 1, 15, -3, 0) op_3955 (v1810[10:0], v2199[13:0], v3955[14:0]); // 3.0
    wire [14:0] v3956; shift_adder #(12, 13, 1, 1, 15, -3, 0) op_3956 (v2200[11:0], v792[12:0], v3956[14:0]); // 3.0
    wire [15:0] v3957; shift_adder #(15, 11, 1, 1, 16, 4, 0) op_3957 (v2201[14:0], v2202[10:0], v3957[15:0]); // 3.0
    wire [26:0] v3958; shift_adder #(11, 26, 1, 1, 27, -16, 0) op_3958 (v2194[10:0], v2203[25:0], v3958[26:0]); // 3.0
    wire [26:0] v3959; shift_adder #(8, 21, 1, 1, 27, -18, 0) op_3959 (v85[7:0], v2204[20:0], v3959[26:0]); // 3.0
    wire [14:0] v3960; shift_adder #(13, 14, 1, 1, 15, 1, 0) op_3960 (v1459[12:0], v2205[13:0], v3960[14:0]); // 3.0
    wire [21:0] v3961; shift_adder #(21, 14, 1, 1, 22, 7, 0) op_3961 (v2206[20:0], v2207[13:0], v3961[21:0]); // 3.0
    wire [19:0] v3962; shift_adder #(13, 18, 1, 1, 20, 2, 1) op_3962 (v524[12:0], v2208[17:0], v3962[19:0]); // 3.0
    wire [15:0] v3963; shift_adder #(16, 14, 1, 1, 16, 1, 0) op_3963 (v2209[15:0], v2147[13:0], v3963[15:0]); // 3.0
    wire [12:0] v3964; shift_adder #(12, 12, 1, 1, 13, 0, 0) op_3964 (v863[11:0], v1893[11:0], v3964[12:0]); // 3.0
    wire [15:0] v3965; shift_adder #(13, 14, 1, 1, 16, -3, 0) op_3965 (v845[12:0], v2210[13:0], v3965[15:0]); // 3.0
    wire [21:0] v3966; shift_adder #(13, 12, 1, 1, 22, -9, 1) op_3966 (v506[12:0], v1745[11:0], v3966[21:0]); // 3.0
    wire [14:0] v3967; shift_adder #(11, 14, 1, 1, 15, 1, 0) op_3967 (v255[10:0], v2075[13:0], v3967[14:0]); // 3.0
    wire [21:0] v3968; shift_adder #(20, 21, 1, 1, 22, -1, 0) op_3968 (v1824[19:0], v1788[20:0], v3968[21:0]); // 3.0
    wire [23:0] v3969; shift_adder #(16, 21, 1, 1, 24, -8, 0) op_3969 (v2211[15:0], v2212[20:0], v3969[23:0]); // 3.0
    wire [23:0] v3970; shift_adder #(16, 23, 1, 1, 24, -8, 0) op_3970 (v1238[15:0], v1733[22:0], v3970[23:0]); // 3.0
    wire [14:0] v3971; shift_adder #(12, 13, 1, 1, 15, -3, 0) op_3971 (v2213[11:0], v2214[12:0], v3971[14:0]); // 3.0
    wire [18:0] v3972; shift_adder #(13, 18, 1, 1, 19, -6, 0) op_3972 (v2215[12:0], v2216[17:0], v3972[18:0]); // 3.0
    wire [16:0] v3973; shift_adder #(16, 12, 1, 1, 17, 4, 0) op_3973 (v1091[15:0], v2116[11:0], v3973[16:0]); // 3.0
    wire [14:0] v3974; shift_adder #(14, 15, 1, 1, 15, 0, 0) op_3974 (v2217[13:0], v1629[14:0], v3974[14:0]); // 3.0
    wire [13:0] v3975; shift_adder #(13, 12, 1, 1, 14, 1, 0) op_3975 (v2218[12:0], v2219[11:0], v3975[13:0]); // 3.0
    wire [24:0] v3976; shift_adder #(14, 25, 1, 1, 25, -9, 0) op_3976 (v975[13:0], v2220[24:0], v3976[24:0]); // 3.0
    wire [15:0] v3977; shift_adder #(14, 11, 1, 1, 16, 4, 0) op_3977 (v1818[13:0], v1054[10:0], v3977[15:0]); // 3.0
    wire [15:0] v3978; shift_adder #(15, 13, 1, 1, 16, 2, 0) op_3978 (v2221[14:0], v1621[12:0], v3978[15:0]); // 3.0
    wire [23:0] v3979; shift_adder #(11, 21, 1, 1, 24, 3, 0) op_3979 (v215[10:0], v1168[20:0], v3979[23:0]); // 3.0
    wire [14:0] v3980; shift_adder #(14, 14, 1, 1, 15, 0, 0) op_3980 (v2222[13:0], v2223[13:0], v3980[14:0]); // 3.0
    wire [17:0] v3981; shift_adder #(17, 16, 1, 1, 18, 2, 0) op_3981 (v2224[16:0], v849[15:0], v3981[17:0]); // 3.0
    wire [14:0] v3982; shift_adder #(14, 12, 1, 1, 15, 2, 0) op_3982 (v1317[13:0], v1283[11:0], v3982[14:0]); // 3.0
    wire [25:0] v3983; shift_adder #(9, 13, 1, 1, 26, -16, 0) op_3983 (v637[8:0], v2225[12:0], v3983[25:0]); // 3.0
    wire [18:0] v3984; shift_adder #(17, 13, 1, 1, 19, 5, 0) op_3984 (v2226[16:0], v1588[12:0], v3984[18:0]); // 3.0
    wire [22:0] v3985; shift_adder #(12, 22, 1, 1, 23, -9, 0) op_3985 (v2227[11:0], v1345[21:0], v3985[22:0]); // 3.0
    wire [30:0] v3986; shift_adder #(30, 12, 1, 1, 31, 18, 0) op_3986 (v2228[29:0], v2229[11:0], v3986[30:0]); // 3.0
    wire [26:0] v3987; shift_adder #(26, 22, 1, 1, 27, 4, 0) op_3987 (v1751[25:0], v1355[21:0], v3987[26:0]); // 3.0
    wire [18:0] v3988; shift_adder #(11, 15, 1, 1, 19, -8, 1) op_3988 (v250[10:0], v1858[14:0], v3988[18:0]); // 3.0
    wire [34:0] v3989; shift_adder #(13, 33, 1, 1, 35, -21, 0) op_3989 (v2225[12:0], v1953[32:0], v3989[34:0]); // 3.0
    wire [24:0] v3990; shift_adder #(23, 18, 1, 1, 25, -2, 1) op_3990 (v2114[22:0], v2230[17:0], v3990[24:0]); // 3.0
    wire [35:0] v3991; shift_adder #(12, 10, 1, 1, 36, 26, 1) op_3991 (v2231[11:0], v705[9:0], v3991[35:0]); // 3.0
    wire [16:0] v3992; shift_adder #(15, 12, 1, 1, 17, 4, 0) op_3992 (v2232[14:0], v2233[11:0], v3992[16:0]); // 3.0
    wire [12:0] v3993; shift_adder #(11, 13, 1, 1, 13, 0, 0) op_3993 (v135[10:0], v2065[12:0], v3993[12:0]); // 3.0
    wire [13:0] v3994; shift_adder #(11, 13, 1, 1, 14, -2, 0) op_3994 (v2234[10:0], v2235[12:0], v3994[13:0]); // 3.0
    wire [13:0] v3995; shift_adder #(13, 13, 1, 1, 14, 0, 0) op_3995 (v2236[12:0], v1209[12:0], v3995[13:0]); // 3.0
    wire [31:0] v3996; shift_adder #(11, 14, 1, 1, 32, 18, 0) op_3996 (v209[10:0], v1834[13:0], v3996[31:0]); // 3.0
    wire [31:0] v3997; shift_adder #(8, 12, 1, 1, 32, 20, 1) op_3997 (v69[7:0], v1977[11:0], v3997[31:0]); // 3.0
    wire [16:0] v3998; shift_adder #(15, 13, 1, 1, 17, 3, 0) op_3998 (v2237[14:0], v1696[12:0], v3998[16:0]); // 3.0
    wire [34:0] v3999; shift_adder #(12, 34, 1, 1, 35, -22, 0) op_3999 (v2238[11:0], v2239[33:0], v3999[34:0]); // 3.0
    wire [17:0] v4000; shift_adder #(13, 17, 1, 1, 18, -4, 0) op_4000 (v2218[12:0], v982[16:0], v4000[17:0]); // 3.0
    wire [36:0] v4001; shift_adder #(12, 13, 1, 1, 37, -25, 1) op_4001 (v1512[11:0], v2240[12:0], v4001[36:0]); // 3.0
    wire [12:0] v4002; shift_adder #(11, 13, 1, 1, 13, 0, 0) op_4002 (v2241[10:0], v845[12:0], v4002[12:0]); // 3.0
    wire [18:0] v4003; shift_adder #(11, 13, 1, 1, 19, 6, 1) op_4003 (v323[10:0], v1202[12:0], v4003[18:0]); // 3.0
    wire [21:0] v4004; shift_adder #(12, 21, 1, 1, 22, -9, 0) op_4004 (v825[11:0], v1191[20:0], v4004[21:0]); // 3.0
    wire [14:0] v4005; shift_adder #(15, 12, 1, 1, 15, 0, 0) op_4005 (v1006[14:0], v797[11:0], v4005[14:0]); // 3.0
    wire [16:0] v4006; shift_adder #(16, 14, 1, 1, 17, 3, 0) op_4006 (v1827[15:0], v2242[13:0], v4006[16:0]); // 3.0
    wire [18:0] v4007; shift_adder #(11, 16, 1, 1, 19, 3, 1) op_4007 (v303[10:0], v1899[15:0], v4007[18:0]); // 3.0
    wire [16:0] v4008; shift_adder #(13, 15, 1, 1, 17, -3, 0) op_4008 (v1670[12:0], v2243[14:0], v4008[16:0]); // 3.0
    wire [15:0] v4009; shift_adder #(12, 14, 1, 1, 16, -3, 0) op_4009 (v1147[11:0], v2244[13:0], v4009[15:0]); // 3.0
    wire [13:0] v4010; shift_adder #(13, 13, 1, 1, 14, -1, 0) op_4010 (v882[12:0], v932[12:0], v4010[13:0]); // 3.0
    wire [14:0] v4011; shift_adder #(12, 13, 1, 1, 15, -3, 0) op_4011 (v2245[11:0], v1819[12:0], v4011[14:0]); // 3.0
    wire [16:0] v4012; shift_adder #(12, 16, 1, 1, 17, -4, 0) op_4012 (v1077[11:0], v2246[15:0], v4012[16:0]); // 3.0
    wire [16:0] v4013; shift_adder #(16, 12, 1, 1, 17, 4, 0) op_4013 (v1201[15:0], v1726[11:0], v4013[16:0]); // 3.0
    wire [15:0] v4014; shift_adder #(13, 14, 1, 1, 16, -2, 0) op_4014 (v2170[12:0], v2134[13:0], v4014[15:0]); // 3.0
    wire [23:0] v4015; shift_adder #(15, 23, 1, 1, 24, -9, 0) op_4015 (v2044[14:0], v1842[22:0], v4015[23:0]); // 3.0
    wire [19:0] v4016; shift_adder #(19, 11, 1, 1, 20, 7, 0) op_4016 (v2052[18:0], v1358[10:0], v4016[19:0]); // 3.0
    wire [14:0] v4017; shift_adder #(12, 13, 1, 1, 15, -2, 0) op_4017 (v1862[11:0], v1295[12:0], v4017[14:0]); // 3.0
    wire [18:0] v4018; shift_adder #(18, 14, 1, 1, 19, 4, 0) op_4018 (v2208[17:0], v2091[13:0], v4018[18:0]); // 3.0
    wire [16:0] v4019; shift_adder #(16, 12, 1, 1, 17, 3, 0) op_4019 (v1389[15:0], v2247[11:0], v4019[16:0]); // 3.0
    wire [17:0] v4020; shift_adder #(14, 17, 1, 1, 18, -4, 1) op_4020 (v1250[13:0], v890[16:0], v4020[17:0]); // 3.0
    wire [14:0] v4021; shift_adder #(12, 13, 1, 1, 15, -2, 0) op_4021 (v2017[11:0], v1070[12:0], v4021[14:0]); // 3.0
    wire [19:0] v4022; shift_adder #(15, 13, 1, 1, 20, 7, 0) op_4022 (v471[14:0], v1736[12:0], v4022[19:0]); // 3.0
    wire [17:0] v4023; shift_adder #(10, 12, 1, 1, 18, -8, 1) op_4023 (v463[9:0], v1584[11:0], v4023[17:0]); // 3.0
    wire [19:0] v4024; shift_adder #(18, 18, 1, 1, 20, -1, 0) op_4024 (v2248[17:0], v2249[17:0], v4024[19:0]); // 3.0
    wire [22:0] v4025; shift_adder #(21, 12, 1, 1, 23, 11, 0) op_4025 (v994[20:0], v2250[11:0], v4025[22:0]); // 3.0
    wire [13:0] v4026; shift_adder #(12, 12, 1, 1, 14, 1, 0) op_4026 (v2251[11:0], v2252[11:0], v4026[13:0]); // 3.0
    wire [15:0] v4027; shift_adder #(13, 16, 1, 1, 16, 0, 0) op_4027 (v1533[12:0], v2253[15:0], v4027[15:0]); // 3.0
    wire [13:0] v4028; shift_adder #(12, 12, 1, 1, 14, 2, 0) op_4028 (v321[11:0], v873[11:0], v4028[13:0]); // 3.0
    wire [25:0] v4029; shift_adder #(26, 12, 1, 1, 26, 13, 0) op_4029 (v1483[25:0], v1255[11:0], v4029[25:0]); // 3.0
    wire [23:0] v4030; shift_adder #(11, 23, 1, 1, 24, -12, 0) op_4030 (v855[10:0], v2114[22:0], v4030[23:0]); // 3.0
    wire [12:0] v4031; shift_adder #(13, 12, 1, 1, 13, 0, 0) op_4031 (v1783[12:0], v2254[11:0], v4031[12:0]); // 3.0
    wire [15:0] v4032; shift_adder #(13, 15, 1, 1, 16, -3, 0) op_4032 (v1209[12:0], v1010[14:0], v4032[15:0]); // 3.0
    wire [21:0] v4033; shift_adder #(20, 12, 1, 1, 22, 9, 0) op_4033 (v2255[19:0], v2256[11:0], v4033[21:0]); // 3.0
    wire [26:0] v4034; shift_adder #(26, 12, 1, 1, 27, 13, 0) op_4034 (v2257[25:0], v1963[11:0], v4034[26:0]); // 3.0
    wire [23:0] v4035; shift_adder #(13, 24, 1, 1, 24, -8, 0) op_4035 (v915[12:0], v1044[23:0], v4035[23:0]); // 3.0
    wire [27:0] v4036; shift_adder #(19, 27, 1, 1, 28, -8, 0) op_4036 (v1942[18:0], v798[26:0], v4036[27:0]); // 3.0
    wire [15:0] v4037; shift_adder #(14, 15, 1, 1, 16, -1, 0) op_4037 (v1679[13:0], v1833[14:0], v4037[15:0]); // 3.0
    wire [24:0] v4038; shift_adder #(15, 24, 1, 1, 25, -8, 0) op_4038 (v1947[14:0], v1087[23:0], v4038[24:0]); // 3.0
    wire [29:0] v4039; shift_adder #(11, 13, 1, 1, 30, -19, 0) op_4039 (v165[10:0], v2258[12:0], v4039[29:0]); // 3.0
    wire [17:0] v4040; shift_adder #(12, 15, 1, 1, 18, -6, 1) op_4040 (v159[11:0], v1011[14:0], v4040[17:0]); // 3.0
    wire [36:0] v4041; shift_adder #(12, 11, 1, 1, 37, 26, 1) op_4041 (v1986[11:0], v320[10:0], v4041[36:0]); // 3.0
    wire [37:0] v4042; shift_adder #(14, 13, 1, 1, 38, -24, 1) op_4042 (v1610[13:0], v2259[12:0], v4042[37:0]); // 3.0
    wire [24:0] v4043; shift_adder #(11, 24, 1, 1, 25, -13, 0) op_4043 (v2260[10:0], v2261[23:0], v4043[24:0]); // 3.0
    wire [39:0] v4044; shift_adder #(39, 36, 1, 1, 40, 4, 0) op_4044 (v2262[38:0], v2263[35:0], v4044[39:0]); // 3.0
    wire [15:0] v4045; shift_adder #(14, 15, 1, 1, 16, -1, 0) op_4045 (v1516[13:0], v1964[14:0], v4045[15:0]); // 3.0
    wire [13:0] v4046; shift_adder #(13, 13, 1, 1, 14, -1, 0) op_4046 (v1138[12:0], v985[12:0], v4046[13:0]); // 3.0
    wire [14:0] v4047; shift_adder #(13, 13, 1, 1, 15, -1, 0) op_4047 (v2264[12:0], v1202[12:0], v4047[14:0]); // 3.0
    wire [13:0] v4048; shift_adder #(11, 13, 1, 1, 14, -2, 1) op_4048 (v132[10:0], v1189[12:0], v4048[13:0]); // 3.0
    wire [15:0] v4049; shift_adder #(14, 14, 1, 1, 16, 2, 0) op_4049 (v1117[13:0], v2265[13:0], v4049[15:0]); // 3.0
    wire [16:0] v4050; shift_adder #(12, 16, 1, 1, 17, -4, 0) op_4050 (v1211[11:0], v2266[15:0], v4050[16:0]); // 3.0
    wire [17:0] v4051; shift_adder #(9, 17, 1, 1, 18, -7, 0) op_4051 (v627[8:0], v1220[16:0], v4051[17:0]); // 3.0
    wire [15:0] v4052; shift_adder #(16, 12, 1, 1, 16, 3, 0) op_4052 (v1169[15:0], v1413[11:0], v4052[15:0]); // 3.0
    wire [15:0] v4053; shift_adder #(15, 13, 1, 1, 16, -1, 0) op_4053 (v2267[14:0], v2268[12:0], v4053[15:0]); // 3.0
    wire [16:0] v4054; shift_adder #(16, 13, 1, 1, 17, 3, 0) op_4054 (v2269[15:0], v1533[12:0], v4054[16:0]); // 3.0
    wire [17:0] v4055; shift_adder #(16, 16, 1, 1, 18, -2, 0) op_4055 (v2270[15:0], v2271[15:0], v4055[17:0]); // 3.0
    wire [30:0] v4056; shift_adder #(30, 14, 1, 1, 31, 16, 0) op_4056 (v2272[29:0], v2273[13:0], v4056[30:0]); // 3.0
    wire [33:0] v4057; shift_adder #(14, 33, 1, 1, 34, -19, 0) op_4057 (v1013[13:0], v1773[32:0], v4057[33:0]); // 3.0
    wire [23:0] v4058; shift_adder #(9, 15, 1, 1, 24, -14, 1) op_4058 (v433[8:0], v815[14:0], v4058[23:0]); // 3.0
    wire [16:0] v4059; shift_adder #(16, 12, 1, 1, 17, 5, 0) op_4059 (v1152[15:0], v2274[11:0], v4059[16:0]); // 3.0
    wire [14:0] v4060; shift_adder #(14, 13, 1, 1, 15, 1, 0) op_4060 (v2275[13:0], v1294[12:0], v4060[14:0]); // 3.0
    wire [31:0] v4061; shift_adder #(19, 32, 1, 1, 32, -11, 0) op_4061 (v1748[18:0], v1318[31:0], v4061[31:0]); // 3.0
    wire [15:0] v4062; shift_adder #(14, 14, 1, 1, 16, -1, 0) op_4062 (v2008[13:0], v2276[13:0], v4062[15:0]); // 3.0
    wire [12:0] v4063; shift_adder #(13, 12, 1, 1, 13, 0, 1) op_4063 (v882[12:0], v279[11:0], v4063[12:0]); // 3.0
    wire [15:0] v4064; shift_adder #(11, 12, 1, 1, 16, -5, 0) op_4064 (v298[10:0], v1498[11:0], v4064[15:0]); // 3.0
    wire [28:0] v4065; shift_adder #(17, 28, 1, 1, 29, -12, 0) op_4065 (v2277[16:0], v2029[27:0], v4065[28:0]); // 3.0
    wire [27:0] v4066; shift_adder #(12, 27, 1, 1, 28, -15, 0) op_4066 (v1555[11:0], v1271[26:0], v4066[27:0]); // 3.0
    wire [27:0] v4067; shift_adder #(27, 15, 1, 1, 28, 12, 0) op_4067 (v2278[26:0], v1690[14:0], v4067[27:0]); // 3.0
    wire [22:0] v4068; shift_adder #(17, 21, 1, 1, 23, -5, 0) op_4068 (v783[16:0], v2279[20:0], v4068[22:0]); // 3.0
    wire [17:0] v4069; shift_adder #(17, 13, 1, 1, 18, -1, 0) op_4069 (v2280[16:0], v2281[12:0], v4069[17:0]); // 3.0
    wire [19:0] v4070; shift_adder #(13, 18, 1, 1, 20, -6, 0) op_4070 (v2066[12:0], v1884[17:0], v4070[19:0]); // 3.0
    wire [19:0] v4071; shift_adder #(19, 14, 1, 1, 20, 5, 0) op_4071 (v782[18:0], v2282[13:0], v4071[19:0]); // 3.0
    wire [13:0] v4072; shift_adder #(12, 13, 1, 1, 14, -1, 0) op_4072 (v2283[11:0], v826[12:0], v4072[13:0]); // 3.0
    wire [14:0] v4073; shift_adder #(13, 13, 1, 1, 15, -1, 0) op_4073 (v996[12:0], v2284[12:0], v4073[14:0]); // 3.0
    wire [12:0] v4074; shift_adder #(10, 13, 1, 1, 13, -1, 1) op_4074 (v549[9:0], v1433[12:0], v4074[12:0]); // 3.0
    wire [13:0] v4075; shift_adder #(13, 12, 1, 1, 14, 1, 0) op_4075 (v2285[12:0], v2286[11:0], v4075[13:0]); // 3.0
    wire [16:0] v4076; shift_adder #(14, 16, 1, 1, 17, 1, 0) op_4076 (v1817[13:0], v970[15:0], v4076[16:0]); // 3.0
    wire [13:0] v4077; shift_adder #(13, 12, 1, 1, 14, 1, 0) op_4077 (v790[12:0], v2238[11:0], v4077[13:0]); // 3.0
    wire [14:0] v4078; shift_adder #(11, 15, 1, 1, 15, -3, 0) op_4078 (v233[10:0], v1027[14:0], v4078[14:0]); // 3.0
    wire [20:0] v4079; shift_adder #(14, 21, 1, 1, 21, -5, 0) op_4079 (v899[13:0], v1586[20:0], v4079[20:0]); // 3.0
    wire [14:0] v4080; shift_adder #(14, 12, 1, 1, 15, 3, 0) op_4080 (v2287[13:0], v929[11:0], v4080[14:0]); // 3.0
    wire [17:0] v4081; shift_adder #(13, 15, 1, 1, 18, -5, 0) op_4081 (v1279[12:0], v2068[14:0], v4081[17:0]); // 3.0
    wire [18:0] v4082; shift_adder #(14, 18, 1, 1, 19, -4, 0) op_4082 (v2288[13:0], v2289[17:0], v4082[18:0]); // 3.0
    wire [17:0] v4083; shift_adder #(17, 15, 1, 1, 18, -1, 0) op_4083 (v1118[16:0], v2068[14:0], v4083[17:0]); // 3.0
    wire [31:0] v4084; shift_adder #(10, 32, 1, 1, 32, -20, 0) op_4084 (v2290[9:0], v2291[31:0], v4084[31:0]); // 3.0
    wire [13:0] v4085; shift_adder #(12, 12, 1, 1, 14, -1, 0) op_4085 (v2292[11:0], v2071[11:0], v4085[13:0]); // 3.0
    wire [13:0] v4086; shift_adder #(13, 11, 1, 1, 14, 2, 0) op_4086 (v1295[12:0], v2293[10:0], v4086[13:0]); // 3.0
    wire [13:0] v4087; shift_adder #(12, 13, 1, 1, 14, -1, 0) op_4087 (v2294[11:0], v2295[12:0], v4087[13:0]); // 3.0
    wire [24:0] v4088; shift_adder #(15, 24, 1, 1, 25, -9, 0) op_4088 (v1265[14:0], v2181[23:0], v4088[24:0]); // 3.0
    wire [28:0] v4089; shift_adder #(10, 21, 1, 1, 29, -19, 1) op_4089 (v291[9:0], v2296[20:0], v4089[28:0]); // 3.0
    wire [16:0] v4090; shift_adder #(17, 12, 1, 1, 17, 2, 0) op_4090 (v2297[16:0], v1641[11:0], v4090[16:0]); // 3.0
    wire [22:0] v4091; shift_adder #(13, 22, 1, 1, 23, -8, 0) op_4091 (v2298[12:0], v1562[21:0], v4091[22:0]); // 3.0
    wire [25:0] v4092; shift_adder #(17, 26, 1, 1, 26, -6, 0) op_4092 (v1674[16:0], v2103[25:0], v4092[25:0]); // 3.0
    wire [32:0] v4093; shift_adder #(18, 32, 1, 1, 33, -15, 0) op_4093 (v2299[17:0], v2291[31:0], v4093[32:0]); // 3.0
    wire [26:0] v4094; shift_adder #(27, 17, 1, 1, 27, 9, 0) op_4094 (v2300[26:0], v2301[16:0], v4094[26:0]); // 3.0
    wire [34:0] v4095; shift_adder #(12, 10, 1, 1, 35, 25, 1) op_4095 (v2302[11:0], v722[9:0], v4095[34:0]); // 3.0
    wire [15:0] v4096; shift_adder #(15, 12, 1, 1, 16, 3, 0) op_4096 (v1417[14:0], v2303[11:0], v4096[15:0]); // 3.0
    wire [36:0] v4097; shift_adder #(12, 12, 1, 1, 37, -25, 1) op_4097 (v2305[11:0], v1730[11:0], v4097[36:0]); // 3.0
    wire [13:0] v4098; shift_adder #(12, 13, 1, 1, 14, -1, 0) op_4098 (v1147[11:0], v2258[12:0], v4098[13:0]); // 3.0
    wire [16:0] v4099; shift_adder #(14, 16, 1, 1, 17, -2, 0) op_4099 (v1507[13:0], v2088[15:0], v4099[16:0]); // 3.0
    wire [14:0] v4100; shift_adder #(11, 14, 1, 1, 15, -3, 0) op_4100 (v1273[10:0], v1007[13:0], v4100[14:0]); // 3.0
    wire [15:0] v4101; shift_adder #(15, 13, 1, 1, 16, 2, 0) op_4101 (v1867[14:0], v2306[12:0], v4101[15:0]); // 3.0
    wire [12:0] v4102; shift_adder #(12, 12, 1, 1, 13, 1, 0) op_4102 (v1534[11:0], v2019[11:0], v4102[12:0]); // 3.0
    wire [35:0] v4103; shift_adder #(35, 34, 1, 1, 36, 1, 0) op_4103 (v2307[34:0], v2308[33:0], v4103[35:0]); // 3.0
    wire [18:0] v4104; shift_adder #(19, 14, 1, 1, 19, 3, 0) op_4104 (v1701[18:0], v2309[13:0], v4104[18:0]); // 3.0
    wire [16:0] v4105; shift_adder #(17, 14, 1, 1, 17, 1, 0) op_4105 (v1485[16:0], v1039[13:0], v4105[16:0]); // 3.0
    wire [15:0] v4106; shift_adder #(15, 13, 1, 1, 16, 1, 0) op_4106 (v1387[14:0], v2310[12:0], v4106[15:0]); // 3.0
    wire [29:0] v4107; shift_adder #(24, 28, 1, 1, 30, -6, 0) op_4107 (v1622[23:0], v2311[27:0], v4107[29:0]); // 3.0
    wire [15:0] v4108; shift_adder #(15, 15, 1, 1, 16, 0, 0) op_4108 (v886[14:0], v1285[14:0], v4108[15:0]); // 3.0
    wire [25:0] v4109; shift_adder #(26, 24, 1, 1, 26, 1, 0) op_4109 (v2312[25:0], v2261[23:0], v4109[25:0]); // 3.0
    wire [24:0] v4110; shift_adder #(12, 24, 1, 1, 25, -12, 0) op_4110 (v2313[11:0], v1729[23:0], v4110[24:0]); // 3.0
    wire [24:0] v4111; shift_adder #(16, 24, 1, 1, 25, -9, 0) op_4111 (v1541[15:0], v2314[23:0], v4111[24:0]); // 3.0
    wire [13:0] v4112; shift_adder #(13, 12, 1, 1, 14, 1, 0) op_4112 (v1941[12:0], v1370[11:0], v4112[13:0]); // 3.0
    wire [24:0] v4113; shift_adder #(12, 23, 1, 1, 25, -12, 0) op_4113 (v2315[11:0], v1645[22:0], v4113[24:0]); // 3.0
    wire [21:0] v4114; shift_adder #(17, 18, 1, 1, 22, -5, 1) op_4114 (v348[16:0], v2025[17:0], v4114[21:0]); // 3.0
    wire [25:0] v4115; shift_adder #(14, 25, 1, 1, 26, -11, 0) op_4115 (v1509[13:0], v1396[24:0], v4115[25:0]); // 3.0
    wire [13:0] v4116; shift_adder #(12, 12, 1, 1, 14, 1, 1) op_4116 (v387[11:0], v1399[11:0], v4116[13:0]); // 3.0
    wire [14:0] v4117; shift_adder #(12, 14, 1, 1, 15, -1, 0) op_4117 (v1498[11:0], v2316[13:0], v4117[14:0]); // 3.0
    wire [23:0] v4118; shift_adder #(18, 22, 1, 1, 24, -6, 0) op_4118 (v949[17:0], v1192[21:0], v4118[23:0]); // 3.0
    wire [21:0] v4119; shift_adder #(21, 20, 1, 1, 22, 1, 0) op_4119 (v1212[20:0], v1983[19:0], v4119[21:0]); // 3.0
    wire [21:0] v4120; shift_adder #(8, 12, 1, 1, 22, 10, 1) op_4120 (v82[7:0], v1077[11:0], v4120[21:0]); // 3.0
    wire [19:0] v4121; shift_adder #(11, 19, 1, 1, 20, -8, 0) op_4121 (v1800[10:0], v2317[18:0], v4121[19:0]); // 3.0
    wire [19:0] v4122; shift_adder #(13, 19, 1, 1, 20, -6, 0) op_4122 (v1078[12:0], v782[18:0], v4122[19:0]); // 3.0
    wire [14:0] v4123; shift_adder #(12, 14, 1, 1, 15, -2, 0) op_4123 (v1558[11:0], v2318[13:0], v4123[14:0]); // 3.0
    wire [17:0] v4124; shift_adder #(13, 17, 1, 1, 18, -4, 0) op_4124 (v1524[12:0], v1540[16:0], v4124[17:0]); // 3.0
    wire [19:0] v4125; shift_adder #(17, 18, 1, 1, 20, -3, 0) op_4125 (v1236[16:0], v1851[17:0], v4125[19:0]); // 3.0
    wire [12:0] v4126; shift_adder #(12, 13, 1, 1, 13, 0, 0) op_4126 (v825[11:0], v1326[12:0], v4126[12:0]); // 3.0
    wire [17:0] v4127; shift_adder #(12, 18, 1, 1, 18, -4, 0) op_4127 (v1278[11:0], v2319[17:0], v4127[17:0]); // 3.0
    wire [15:0] v4128; shift_adder #(16, 12, 1, 1, 16, 3, 0) op_4128 (v2320[15:0], v879[11:0], v4128[15:0]); // 3.0
    wire [16:0] v4129; shift_adder #(14, 16, 1, 1, 17, 1, 0) op_4129 (v950[13:0], v946[15:0], v4129[16:0]); // 3.0
    wire [14:0] v4130; shift_adder #(11, 14, 1, 1, 15, -3, 0) op_4130 (v2321[10:0], v1522[13:0], v4130[14:0]); // 3.0
    wire [19:0] v4131; shift_adder #(19, 12, 1, 1, 20, 7, 0) op_4131 (v2322[18:0], v1493[11:0], v4131[19:0]); // 3.0
    wire [17:0] v4132; shift_adder #(15, 18, 1, 1, 18, -2, 0) op_4132 (v2323[14:0], v2324[17:0], v4132[17:0]); // 3.0
    wire [16:0] v4133; shift_adder #(12, 12, 1, 1, 17, 5, 0) op_4133 (v404[11:0], v2135[11:0], v4133[16:0]); // 3.0
    wire [22:0] v4134; shift_adder #(21, 20, 1, 1, 23, 2, 0) op_4134 (v2279[20:0], v2172[19:0], v4134[22:0]); // 3.0
    wire [18:0] v4135; shift_adder #(12, 18, 1, 1, 19, -6, 0) op_4135 (v1836[11:0], v2325[17:0], v4135[18:0]); // 3.0
    wire [22:0] v4136; shift_adder #(22, 13, 1, 1, 23, 9, 0) op_4136 (v2326[21:0], v826[12:0], v4136[22:0]); // 3.0
    wire [16:0] v4137; shift_adder #(14, 16, 1, 1, 17, -2, 0) op_4137 (v2327[13:0], v1414[15:0], v4137[16:0]); // 3.0
    wire [31:0] v4138; shift_adder #(12, 31, 1, 1, 32, -19, 1) op_4138 (v1379[11:0], v641[30:0], v4138[31:0]); // 3.0
    wire [19:0] v4139; shift_adder #(18, 17, 1, 1, 20, 3, 0) op_4139 (v1073[17:0], v2328[16:0], v4139[19:0]); // 3.0
    wire [32:0] v4140; shift_adder #(28, 33, 1, 1, 33, -2, 0) op_4140 (v2311[27:0], v2329[32:0], v4140[32:0]); // 3.0
    wire [13:0] v4141; shift_adder #(12, 12, 1, 1, 14, -1, 0) op_4141 (v2124[11:0], v2330[11:0], v4141[13:0]); // 3.0
    wire [23:0] v4142; shift_adder #(23, 19, 1, 1, 24, 5, 0) op_4142 (v1141[22:0], v1210[18:0], v4142[23:0]); // 3.0
    wire [37:0] v4143; shift_adder #(14, 38, 1, 1, 38, -23, 0) op_4143 (v2331[13:0], v2332[37:0], v4143[37:0]); // 3.0
    wire [13:0] v4144; shift_adder #(13, 12, 1, 1, 14, -1, 0) op_4144 (v2333[12:0], v2334[11:0], v4144[13:0]); // 3.0
    wire [12:0] v4145; shift_adder #(11, 12, 1, 1, 13, -1, 0) op_4145 (v2335[10:0], v1069[11:0], v4145[12:0]); // 3.0
    wire [14:0] v4146; shift_adder #(15, 13, 1, 1, 15, 0, 0) op_4146 (v2336[14:0], v1375[12:0], v4146[14:0]); // 3.0
    wire [18:0] v4147; shift_adder #(19, 13, 1, 1, 19, 1, 0) op_4147 (v1945[18:0], v1422[12:0], v4147[18:0]); // 3.0
    wire [18:0] v4148; shift_adder #(12, 18, 1, 1, 19, -5, 0) op_4148 (v1655[11:0], v853[17:0], v4148[18:0]); // 3.0
    wire [13:0] v4149; shift_adder #(13, 13, 1, 1, 14, 0, 0) op_4149 (v1336[12:0], v1741[12:0], v4149[13:0]); // 3.0
    wire [12:0] v4150; shift_adder #(12, 12, 1, 1, 13, 0, 0) op_4150 (v2337[11:0], v1726[11:0], v4150[12:0]); // 3.0
    wire [13:0] v4151; shift_adder #(12, 12, 1, 1, 14, -1, 0) op_4151 (v1888[11:0], v2338[11:0], v4151[13:0]); // 3.0
    wire [13:0] v4152; shift_adder #(10, 12, 1, 1, 14, -3, 0) op_4152 (v2339[9:0], v2340[11:0], v4152[13:0]); // 3.0
    wire [19:0] v4153; shift_adder #(19, 12, 1, 1, 20, 7, 0) op_4153 (v1321[18:0], v2341[11:0], v4153[19:0]); // 3.0
    wire [39:0] v4154; shift_adder #(33, 39, 1, 1, 40, -5, 0) op_4154 (v1441[32:0], v2342[38:0], v4154[39:0]); // 3.0
    wire [13:0] v4155; shift_adder #(13, 12, 1, 1, 14, 1, 0) op_4155 (v1569[12:0], v1082[11:0], v4155[13:0]); // 3.0
    wire [16:0] v4156; shift_adder #(17, 13, 1, 1, 17, 2, 1) op_4156 (v1175[16:0], v1438[12:0], v4156[16:0]); // 3.0
    wire [29:0] v4157; shift_adder #(28, 30, 1, 1, 30, -1, 0) op_4157 (v1528[27:0], v2343[29:0], v4157[29:0]); // 3.0
    wire [19:0] v4158; shift_adder #(19, 19, 1, 1, 20, -1, 0) op_4158 (v1814[18:0], v2197[18:0], v4158[19:0]); // 3.0
    wire [26:0] v4159; shift_adder #(20, 26, 1, 1, 27, -5, 0) op_4159 (v1603[19:0], v2344[25:0], v4159[26:0]); // 3.0
    wire [25:0] v4160; shift_adder #(9, 15, 1, 1, 26, -17, 1) op_4160 (v351[8:0], v1721[14:0], v4160[25:0]); // 3.0
    wire [30:0] v4161; shift_adder #(31, 17, 1, 1, 31, 12, 0) op_4161 (v1693[30:0], v2345[16:0], v4161[30:0]); // 3.0
    wire [14:0] v4162; shift_adder #(11, 13, 1, 1, 15, -4, 0) op_4162 (v2346[10:0], v932[12:0], v4162[14:0]); // 3.0
    wire [14:0] v4163; shift_adder #(14, 12, 1, 1, 15, 1, 0) op_4163 (v2199[13:0], v1171[11:0], v4163[14:0]); // 3.0
    wire [24:0] v4164; shift_adder #(8, 13, 1, 1, 25, -16, 0) op_4164 (v121[7:0], v985[12:0], v4164[24:0]); // 3.0
    wire [25:0] v4165; shift_adder #(12, 26, 1, 1, 26, -10, 0) op_4165 (v512[11:0], v2347[25:0], v4165[25:0]); // 3.0
    wire [17:0] v4166; shift_adder #(12, 18, 1, 1, 18, -4, 0) op_4166 (v1190[11:0], v872[17:0], v4166[17:0]); // 3.0
    wire [16:0] v4167; shift_adder #(12, 14, 1, 1, 17, -4, 0) op_4167 (v2348[11:0], v2134[13:0], v4167[16:0]); // 3.0
    wire [25:0] v4168; shift_adder #(25, 22, 1, 1, 26, 4, 1) op_4168 (v537[24:0], v2349[21:0], v4168[25:0]); // 3.0
    wire [21:0] v4169; shift_adder #(13, 20, 1, 1, 22, -8, 0) op_4169 (v2350[12:0], v2351[19:0], v4169[21:0]); // 3.0
    wire [17:0] v4170; shift_adder #(16, 14, 1, 1, 18, 3, 0) op_4170 (v927[15:0], v1859[13:0], v4170[17:0]); // 3.0
    wire [15:0] v4171; shift_adder #(13, 14, 1, 1, 16, -2, 0) op_4171 (v1074[12:0], v899[13:0], v4171[15:0]); // 3.0
    wire [20:0] v4172; shift_adder #(12, 20, 1, 1, 21, -7, 0) op_4172 (v2352[11:0], v1289[19:0], v4172[20:0]); // 3.0
    wire [13:0] v4173; shift_adder #(13, 13, 1, 1, 14, 0, 0) op_4173 (v2353[12:0], v2354[12:0], v4173[13:0]); // 3.0
    wire [13:0] v4174; shift_adder #(11, 13, 1, 1, 14, -2, 0) op_4174 (v1284[10:0], v1949[12:0], v4174[13:0]); // 3.0
    wire [23:0] v4175; shift_adder #(15, 22, 1, 1, 24, -9, 0) op_4175 (v2267[14:0], v2032[21:0], v4175[23:0]); // 3.0
    wire [21:0] v4176; shift_adder #(16, 22, 1, 1, 22, -5, 0) op_4176 (v1382[15:0], v2355[21:0], v4176[21:0]); // 3.0
    wire [13:0] v4177; shift_adder #(11, 11, 1, 1, 14, 2, 1) op_4177 (v374[10:0], v785[10:0], v4177[13:0]); // 3.0
    wire [27:0] v4178; shift_adder #(27, 14, 1, 1, 28, 14, 0) op_4178 (v1989[26:0], v2356[13:0], v4178[27:0]); // 3.0
    wire [21:0] v4179; shift_adder #(11, 21, 1, 1, 22, 1, 0) op_4179 (v338[10:0], v1266[20:0], v4179[21:0]); // 3.0
    wire [15:0] v4180; shift_adder #(14, 15, 1, 1, 16, -1, 0) op_4180 (v1126[13:0], v2357[14:0], v4180[15:0]); // 3.0
    wire [18:0] v4181; shift_adder #(14, 17, 1, 1, 19, -4, 0) op_4181 (v2273[13:0], v1392[16:0], v4181[18:0]); // 3.0
    wire [23:0] v4182; shift_adder #(13, 24, 1, 1, 24, -10, 0) op_4182 (v2358[12:0], v1515[23:0], v4182[23:0]); // 3.0
    wire [27:0] v4183; shift_adder #(27, 18, 1, 1, 28, 9, 0) op_4183 (v2359[26:0], v2360[17:0], v4183[27:0]); // 3.0
    wire [13:0] v4184; shift_adder #(13, 11, 1, 1, 14, 1, 0) op_4184 (v1324[12:0], v1943[10:0], v4184[13:0]); // 3.0
    wire [26:0] v4185; shift_adder #(25, 26, 1, 1, 27, 1, 0) op_4185 (v2361[24:0], v802[25:0], v4185[26:0]); // 3.0
    wire [16:0] v4186; shift_adder #(16, 16, 1, 1, 17, -1, 0) op_4186 (v1275[15:0], v2362[15:0], v4186[16:0]); // 3.0
    wire [13:0] v4187; shift_adder #(8, 13, 1, 1, 14, -5, 1) op_4187 (v80[7:0], v2298[12:0], v4187[13:0]); // 3.0
    wire [14:0] v4188; shift_adder #(13, 13, 1, 1, 15, 1, 0) op_4188 (v828[12:0], v1074[12:0], v4188[14:0]); // 3.0
    wire [16:0] v4189; shift_adder #(14, 17, 1, 1, 17, -2, 0) op_4189 (v2363[13:0], v1809[16:0], v4189[16:0]); // 3.0
    wire [31:0] v4190; shift_adder #(16, 32, 1, 1, 32, -14, 0) op_4190 (v1606[15:0], v1654[31:0], v4190[31:0]); // 3.0
    wire [17:0] v4191; shift_adder #(17, 13, 1, 1, 18, 3, 0) op_4191 (v1291[16:0], v2031[12:0], v4191[17:0]); // 3.0
    wire [15:0] v4192; shift_adder #(14, 14, 1, 1, 16, -2, 0) op_4192 (v2364[13:0], v1545[13:0], v4192[15:0]); // 3.0
    wire [34:0] v4193; shift_adder #(33, 18, 1, 1, 35, 17, 0) op_4193 (v2365[32:0], v1592[17:0], v4193[34:0]); // 3.0
    wire [18:0] v4194; shift_adder #(13, 19, 1, 1, 19, -5, 0) op_4194 (v793[12:0], v2366[18:0], v4194[18:0]); // 3.0
    wire [14:0] v4195; shift_adder #(14, 10, 1, 1, 15, 4, 0) op_4195 (v2186[13:0], v2104[9:0], v4195[14:0]); // 3.0
    wire [18:0] v4196; shift_adder #(12, 17, 1, 1, 19, -6, 0) op_4196 (v956[11:0], v1519[16:0], v4196[18:0]); // 3.0
    wire [15:0] v4197; shift_adder #(15, 12, 1, 1, 16, 3, 0) op_4197 (v1572[14:0], v2367[11:0], v4197[15:0]); // 3.0
    wire [32:0] v4198; shift_adder #(12, 31, 1, 1, 33, -20, 0) op_4198 (v1105[11:0], v1488[30:0], v4198[32:0]); // 3.0
    wire [39:0] v4199; shift_adder #(15, 15, 1, 1, 40, 25, 1) op_4199 (v2368[14:0], v733[14:0], v4199[39:0]); // 3.0
    wire [16:0] v4200; shift_adder #(16, 11, 1, 1, 17, 5, 0) op_4200 (v970[15:0], v2123[10:0], v4200[16:0]); // 3.0
    wire [13:0] v4201; shift_adder #(13, 13, 1, 1, 14, 0, 0) op_4201 (v2369[12:0], v1046[12:0], v4201[13:0]); // 3.0
    wire [33:0] v4202; shift_adder #(33, 12, 1, 1, 34, 21, 0) op_4202 (v1060[32:0], v1850[11:0], v4202[33:0]); // 3.0
    wire [37:0] v4203; shift_adder #(18, 13, 1, 1, 38, -20, 1) op_4203 (v1094[17:0], v826[12:0], v4203[37:0]); // 3.0
    wire [13:0] v4204; shift_adder #(12, 13, 1, 1, 14, -1, 0) op_4204 (v1829[11:0], v2370[12:0], v4204[13:0]); // 3.0
    wire [14:0] v4205; shift_adder #(11, 13, 1, 1, 15, -3, 0) op_4205 (v2293[10:0], v2371[12:0], v4205[14:0]); // 3.0
    wire [11:0] v4206; shift_adder #(12, 11, 1, 1, 12, 0, 0) op_4206 (v2372[11:0], v2346[10:0], v4206[11:0]); // 3.0
    wire [15:0] v4207; shift_adder #(15, 13, 1, 1, 16, 2, 0) op_4207 (v1879[14:0], v2353[12:0], v4207[15:0]); // 3.0
    wire [24:0] v4208; shift_adder #(25, 16, 1, 1, 25, 8, 0) op_4208 (v2026[24:0], v970[15:0], v4208[24:0]); // 3.0
    wire [18:0] v4209; shift_adder #(12, 17, 1, 1, 19, -7, 0) op_4209 (v2017[11:0], v1546[16:0], v4209[18:0]); // 3.0
    wire [13:0] v4210; shift_adder #(13, 14, 1, 1, 14, 0, 0) op_4210 (v915[12:0], v975[13:0], v4210[13:0]); // 3.0
    wire [20:0] v4211; shift_adder #(21, 19, 1, 1, 21, 1, 0) op_4211 (v1267[20:0], v2052[18:0], v4211[20:0]); // 3.0
    wire [17:0] v4212; shift_adder #(14, 18, 1, 1, 18, -3, 0) op_4212 (v1817[13:0], v1709[17:0], v4212[17:0]); // 3.0
    wire [18:0] v4213; shift_adder #(13, 17, 1, 1, 19, -6, 0) op_4213 (v2141[12:0], v2224[16:0], v4213[18:0]); // 3.0
    wire [17:0] v4214; shift_adder #(17, 15, 1, 1, 18, 1, 0) op_4214 (v2373[16:0], v1932[14:0], v4214[17:0]); // 3.0
    wire [18:0] v4215; shift_adder #(18, 12, 1, 1, 19, 6, 0) op_4215 (v1453[17:0], v1906[11:0], v4215[18:0]); // 3.0
    wire [12:0] v4216; shift_adder #(12, 10, 1, 1, 13, 2, 0) op_4216 (v2374[11:0], v2183[9:0], v4216[12:0]); // 3.0
    wire [14:0] v4217; shift_adder #(13, 13, 1, 1, 15, -1, 0) op_4217 (v2375[12:0], v1397[12:0], v4217[14:0]); // 3.0
    wire [13:0] v4218; shift_adder #(13, 13, 1, 1, 14, 0, 0) op_4218 (v1560[12:0], v2376[12:0], v4218[13:0]); // 3.0
    wire [13:0] v4219; shift_adder #(12, 12, 1, 1, 14, -1, 0) op_4219 (v2377[11:0], v2378[11:0], v4219[13:0]); // 3.0
    wire [15:0] v4220; shift_adder #(14, 14, 1, 1, 16, 2, 0) op_4220 (v2379[13:0], v1575[13:0], v4220[15:0]); // 3.0
    wire [17:0] v4221; shift_adder #(17, 12, 1, 1, 18, 4, 0) op_4221 (v2380[16:0], v1136[11:0], v4221[17:0]); // 3.0
    wire [18:0] v4222; shift_adder #(15, 15, 1, 1, 19, 4, 0) op_4222 (v1107[14:0], v2381[14:0], v4222[18:0]); // 3.0
    wire [12:0] v4223; shift_adder #(12, 12, 1, 1, 13, 1, 0) op_4223 (v820[11:0], v2382[11:0], v4223[12:0]); // 3.0
    wire [15:0] v4224; shift_adder #(11, 15, 1, 1, 16, -4, 0) op_4224 (v2123[10:0], v2383[14:0], v4224[15:0]); // 3.0
    wire [20:0] v4225; shift_adder #(20, 16, 1, 1, 21, 4, 0) op_4225 (v1567[19:0], v2209[15:0], v4225[20:0]); // 3.0
    wire [20:0] v4226; shift_adder #(19, 20, 1, 1, 21, 1, 0) op_4226 (v1009[18:0], v2384[19:0], v4226[20:0]); // 3.0
    wire [22:0] v4227; shift_adder #(23, 13, 1, 1, 23, 9, 0) op_4227 (v1954[22:0], v1375[12:0], v4227[22:0]); // 3.0
    wire [17:0] v4228; shift_adder #(13, 14, 1, 1, 18, 4, 1) op_4228 (v859[12:0], v1300[13:0], v4228[17:0]); // 3.0
    wire [18:0] v4229; shift_adder #(15, 19, 1, 1, 19, -3, 0) op_4229 (v1632[14:0], v776[18:0], v4229[18:0]); // 3.0
    wire [19:0] v4230; shift_adder #(12, 19, 1, 1, 20, -8, 0) op_4230 (v2385[11:0], v1772[18:0], v4230[19:0]); // 3.0
    wire [17:0] v4231; shift_adder #(13, 15, 1, 1, 18, 3, 0) op_4231 (v2386[12:0], v1611[14:0], v4231[17:0]); // 3.0
    wire [14:0] v4232; shift_adder #(13, 13, 1, 1, 15, 2, 0) op_4232 (v1026[12:0], v1356[12:0], v4232[14:0]); // 3.0
    wire [17:0] v4233; shift_adder #(17, 16, 1, 1, 18, -1, 1) op_4233 (v1118[16:0], v1762[15:0], v4233[17:0]); // 3.0
    wire [13:0] v4234; shift_adder #(10, 13, 1, 1, 14, -2, 0) op_4234 (v2290[9:0], v2100[12:0], v4234[13:0]); // 3.0
    wire [25:0] v4235; shift_adder #(12, 26, 1, 1, 26, -13, 0) op_4235 (v1602[11:0], v1338[25:0], v4235[25:0]); // 3.0
    wire [27:0] v4236; shift_adder #(27, 14, 1, 1, 28, 13, 0) op_4236 (v2278[26:0], v2387[13:0], v4236[27:0]); // 3.0
    wire [22:0] v4237; shift_adder #(14, 23, 1, 1, 23, -1, 1) op_4237 (v412[13:0], v1319[22:0], v4237[22:0]); // 3.0
    wire [15:0] v4238; shift_adder #(12, 14, 1, 1, 16, -3, 0) op_4238 (v2388[11:0], v871[13:0], v4238[15:0]); // 3.0
    wire [16:0] v4239; shift_adder #(16, 15, 1, 1, 17, 2, 0) op_4239 (v1275[15:0], v1010[14:0], v4239[16:0]); // 3.0
    wire [18:0] v4240; shift_adder #(18, 13, 1, 1, 19, 5, 0) op_4240 (v2389[17:0], v2390[12:0], v4240[18:0]); // 3.0
    wire [14:0] v4241; shift_adder #(15, 13, 1, 1, 15, 0, 0) op_4241 (v2391[14:0], v2392[12:0], v4241[14:0]); // 3.0
    wire [15:0] v4242; shift_adder #(11, 15, 1, 1, 16, -4, 0) op_4242 (v1943[10:0], v2117[14:0], v4242[15:0]); // 3.0
    wire [23:0] v4243; shift_adder #(18, 23, 1, 1, 24, -6, 0) op_4243 (v2140[17:0], v1842[22:0], v4243[23:0]); // 3.0
    wire [37:0] v4244; shift_adder #(36, 13, 1, 1, 38, 24, 0) op_4244 (v2394[35:0], v2395[12:0], v4244[37:0]); // 3.0
    wire [27:0] v4245; shift_adder #(27, 14, 1, 1, 28, 13, 0) op_4245 (v1260[26:0], v2143[13:0], v4245[27:0]); // 3.0
    wire [12:0] v4246; shift_adder #(11, 12, 1, 1, 13, -1, 0) op_4246 (v1627[10:0], v1708[11:0], v4246[12:0]); // 3.0
    wire [15:0] v4247; shift_adder #(14, 14, 1, 1, 16, -1, 0) op_4247 (v1332[13:0], v1288[13:0], v4247[15:0]); // 3.0
    wire [14:0] v4248; shift_adder #(11, 13, 1, 1, 15, -3, 0) op_4248 (v2095[10:0], v1041[12:0], v4248[14:0]); // 3.0
    wire [14:0] v4249; shift_adder #(14, 12, 1, 1, 15, -1, 0) op_4249 (v2396[13:0], v1475[11:0], v4249[14:0]); // 3.0
    wire [18:0] v4250; shift_adder #(12, 17, 1, 1, 19, -6, 0) op_4250 (v2286[11:0], v2397[16:0], v4250[18:0]); // 3.0
    wire [32:0] v4251; shift_adder #(22, 32, 1, 1, 33, -10, 0) op_4251 (v1988[21:0], v1815[31:0], v4251[32:0]); // 3.0
    wire [21:0] v4252; shift_adder #(18, 20, 1, 1, 22, -3, 0) op_4252 (v2047[17:0], v2398[19:0], v4252[21:0]); // 3.0
    wire [21:0] v4253; shift_adder #(21, 16, 1, 1, 22, 5, 0) op_4253 (v2296[20:0], v1691[15:0], v4253[21:0]); // 3.0
    wire [15:0] v4254; shift_adder #(15, 12, 1, 1, 16, 3, 0) op_4254 (v2243[14:0], v2399[11:0], v4254[15:0]); // 3.0
    wire [24:0] v4255; shift_adder #(24, 13, 1, 1, 25, 11, 0) op_4255 (v1703[23:0], v2400[12:0], v4255[24:0]); // 3.0
    wire [25:0] v4256; shift_adder #(11, 24, 1, 1, 26, -14, 0) op_4256 (v2401[10:0], v2314[23:0], v4256[25:0]); // 3.0
    wire [25:0] v4257; shift_adder #(25, 15, 1, 1, 26, 11, 0) op_4257 (v796[24:0], v1609[14:0], v4257[25:0]); // 3.0
    wire [18:0] v4258; shift_adder #(12, 18, 1, 1, 19, -7, 0) op_4258 (v2402[11:0], v2145[17:0], v4258[18:0]); // 3.0
    wire [23:0] v4259; shift_adder #(14, 23, 1, 1, 24, -9, 0) op_4259 (v1229[13:0], v2403[22:0], v4259[23:0]); // 3.0
    wire [13:0] v4260; shift_adder #(13, 12, 1, 1, 14, 1, 0) op_4260 (v1458[12:0], v825[11:0], v4260[13:0]); // 3.0
    wire [15:0] v4261; shift_adder #(12, 16, 1, 1, 16, -2, 0) op_4261 (v2404[11:0], v901[15:0], v4261[15:0]); // 3.0
    wire [14:0] v4262; shift_adder #(14, 13, 1, 1, 15, -1, 0) op_4262 (v1575[13:0], v920[12:0], v4262[14:0]); // 3.0
    wire [20:0] v4263; shift_adder #(20, 17, 1, 1, 21, -1, 0) op_4263 (v1666[19:0], v1618[16:0], v4263[20:0]); // 3.0
    wire [21:0] v4264; shift_adder #(22, 12, 1, 1, 22, 8, 0) op_4264 (v2349[21:0], v2405[11:0], v4264[21:0]); // 3.0
    wire [22:0] v4265; shift_adder #(22, 15, 1, 1, 23, 7, 0) op_4265 (v906[21:0], v1536[14:0], v4265[22:0]); // 3.0
    wire [16:0] v4266; shift_adder #(17, 13, 1, 1, 17, 1, 0) op_4266 (v2406[16:0], v2407[12:0], v4266[16:0]); // 3.0
    wire [15:0] v4267; shift_adder #(15, 15, 1, 1, 16, 1, 0) op_4267 (v1038[14:0], v1387[14:0], v4267[15:0]); // 3.0
    wire [20:0] v4268; shift_adder #(20, 15, 1, 1, 21, 6, 0) op_4268 (v2255[19:0], v2022[14:0], v4268[20:0]); // 3.0
    wire [17:0] v4269; shift_adder #(12, 15, 1, 1, 18, -5, 0) op_4269 (v1585[11:0], v2323[14:0], v4269[17:0]); // 3.0
    wire [24:0] v4270; shift_adder #(25, 14, 1, 1, 25, 9, 0) op_4270 (v2408[24:0], v2409[13:0], v4270[24:0]); // 3.0
    wire [29:0] v4271; shift_adder #(15, 30, 1, 1, 30, -11, 0) op_4271 (v2099[14:0], v1232[29:0], v4271[29:0]); // 3.0
    wire [27:0] v4272; shift_adder #(25, 28, 1, 1, 28, -2, 0) op_4272 (v1269[24:0], v1803[27:0], v4272[27:0]); // 3.0
    wire [23:0] v4273; shift_adder #(22, 12, 1, 1, 24, 11, 0) op_4273 (v2023[21:0], v2410[11:0], v4273[23:0]); // 3.0
    wire [27:0] v4274; shift_adder #(27, 11, 1, 1, 28, 16, 0) op_4274 (v1657[26:0], v2411[10:0], v4274[27:0]); // 3.0
    wire [14:0] v4275; shift_adder #(13, 14, 1, 1, 15, 0, 0) op_4275 (v932[12:0], v2412[13:0], v4275[14:0]); // 3.0
    wire [20:0] v4276; shift_adder #(20, 13, 1, 1, 21, 8, 0) op_4276 (v1075[19:0], v920[12:0], v4276[20:0]); // 3.0
    wire [16:0] v4277; shift_adder #(16, 15, 1, 1, 17, 1, 0) op_4277 (v2413[15:0], v2414[14:0], v4277[16:0]); // 3.0
    wire [19:0] v4278; shift_adder #(19, 13, 1, 1, 20, 6, 0) op_4278 (v1764[18:0], v1458[12:0], v4278[19:0]); // 3.0
    wire [15:0] v4279; shift_adder #(14, 12, 1, 1, 16, 3, 0) op_4279 (v1381[13:0], v1105[11:0], v4279[15:0]); // 3.0
    wire [23:0] v4280; shift_adder #(22, 21, 1, 1, 24, 3, 0) op_4280 (v2415[21:0], v1864[20:0], v4280[23:0]); // 3.0
    wire [21:0] v4281; shift_adder #(12, 21, 1, 1, 22, -9, 0) op_4281 (v2416[11:0], v1539[20:0], v4281[21:0]); // 3.0
    wire [16:0] v4282; shift_adder #(11, 15, 1, 1, 17, -5, 0) op_4282 (v1419[10:0], v2046[14:0], v4282[16:0]); // 3.0
    wire [13:0] v4283; shift_adder #(14, 12, 1, 1, 14, 0, 0) op_4283 (v2417[13:0], v2418[11:0], v4283[13:0]); // 3.0
    wire [16:0] v4284; shift_adder #(17, 12, 1, 1, 17, 3, 0) op_4284 (v972[16:0], v1694[11:0], v4284[16:0]); // 3.0
    wire [14:0] v4285; shift_adder #(11, 14, 1, 1, 15, -2, 0) op_4285 (v2346[10:0], v2419[13:0], v4285[14:0]); // 3.0
    wire [18:0] v4286; shift_adder #(18, 16, 1, 1, 19, 2, 0) op_4286 (v1005[17:0], v1889[15:0], v4286[18:0]); // 3.0
    wire [16:0] v4287; shift_adder #(11, 16, 1, 1, 17, -3, 0) op_4287 (v885[10:0], v2420[15:0], v4287[16:0]); // 3.0
    wire [37:0] v4288; shift_adder #(12, 10, 1, 1, 38, 28, 1) op_4288 (v1756[11:0], v450[9:0], v4288[37:0]); // 3.0
    wire [13:0] v4289; shift_adder #(12, 13, 1, 1, 14, 0, 0) op_4289 (v1468[11:0], v2421[12:0], v4289[13:0]); // 3.0
    wire [18:0] v4290; shift_adder #(10, 19, 1, 1, 19, -8, 0) op_4290 (v2104[9:0], v2197[18:0], v4290[18:0]); // 3.0
    wire [14:0] v4291; shift_adder #(12, 13, 1, 1, 15, -2, 0) op_4291 (v2422[11:0], v2423[12:0], v4291[14:0]); // 3.0
    wire [16:0] v4292; shift_adder #(17, 12, 1, 1, 17, 3, 0) op_4292 (v1464[16:0], v2424[11:0], v4292[16:0]); // 3.0
    wire [16:0] v4293; shift_adder #(13, 15, 1, 1, 17, -4, 1) op_4293 (v882[12:0], v1832[14:0], v4293[16:0]); // 3.0
    wire [16:0] v4294; shift_adder #(15, 12, 1, 1, 17, 4, 0) op_4294 (v1879[14:0], v2425[11:0], v4294[16:0]); // 3.0
    wire [41:0] v4295; shift_adder #(11, 40, 1, 1, 42, -30, 0) op_4295 (v2426[10:0], v2427[39:0], v4295[41:0]); // 3.0
    wire [13:0] v4296; shift_adder #(11, 12, 1, 1, 14, -2, 0) op_4296 (v2428[10:0], v1669[11:0], v4296[13:0]); // 3.0
    wire [18:0] v4297; shift_adder #(18, 13, 1, 1, 19, 5, 0) op_4297 (v2025[17:0], v845[12:0], v4297[18:0]); // 3.0
    wire [15:0] v4298; shift_adder #(12, 15, 1, 1, 16, -3, 0) op_4298 (v1100[11:0], v2003[14:0], v4298[15:0]); // 3.0
    wire [14:0] v4299; shift_adder #(13, 13, 1, 1, 15, 1, 0) op_4299 (v1074[12:0], v1336[12:0], v4299[14:0]); // 3.0
    wire [12:0] v4300; shift_adder #(12, 12, 1, 1, 13, -1, 0) op_4300 (v2429[11:0], v862[11:0], v4300[12:0]); // 3.0
    wire [14:0] v4301; shift_adder #(11, 14, 1, 1, 15, -3, 0) op_4301 (v2346[10:0], v2430[13:0], v4301[14:0]); // 3.0
    wire [15:0] v4302; shift_adder #(14, 14, 1, 1, 16, 2, 0) op_4302 (v2118[13:0], v1394[13:0], v4302[15:0]); // 3.0
    wire [11:0] v4303; shift_adder #(11, 11, 1, 1, 12, 0, 0) op_4303 (v2431[10:0], v1517[10:0], v4303[11:0]); // 3.0
    wire [29:0] v4304; shift_adder #(30, 15, 1, 1, 30, 10, 0) op_4304 (v2121[29:0], v1583[14:0], v4304[29:0]); // 3.0
    wire [15:0] v4305; shift_adder #(15, 15, 1, 1, 16, 1, 0) op_4305 (v2432[14:0], v2005[14:0], v4305[15:0]); // 3.0
    wire [17:0] v4306; shift_adder #(17, 14, 1, 1, 18, 3, 0) op_4306 (v852[16:0], v2433[13:0], v4306[17:0]); // 3.0
    wire [27:0] v4307; shift_adder #(27, 20, 1, 1, 28, 6, 0) op_4307 (v1687[26:0], v2351[19:0], v4307[27:0]); // 3.0
    wire [27:0] v4308; shift_adder #(24, 25, 1, 1, 28, -4, 0) op_4308 (v1268[23:0], v2361[24:0], v4308[27:0]); // 3.0
    wire [16:0] v4309; shift_adder #(12, 13, 1, 1, 17, -5, 0) op_4309 (v2434[11:0], v2098[12:0], v4309[16:0]); // 3.0
    wire [18:0] v4310; shift_adder #(17, 18, 1, 1, 19, -1, 0) op_4310 (v2277[16:0], v940[17:0], v4310[18:0]); // 3.0
    wire [28:0] v4311; shift_adder #(13, 13, 1, 1, 29, 16, 0) op_4311 (v1024[12:0], v2268[12:0], v4311[28:0]); // 3.0
    wire [26:0] v4312; shift_adder #(12, 15, 1, 1, 27, -15, 1) op_4312 (v336[11:0], v1352[14:0], v4312[26:0]); // 3.0
    wire [23:0] v4313; shift_adder #(13, 24, 1, 1, 24, -10, 0) op_4313 (v1227[12:0], v2435[23:0], v4313[23:0]); // 3.0
    wire [19:0] v4314; shift_adder #(13, 18, 1, 1, 20, -7, 0) op_4314 (v2421[12:0], v977[17:0], v4314[19:0]); // 3.0
    wire [12:0] v4315; shift_adder #(12, 9, 1, 1, 13, 3, 1) op_4315 (v825[11:0], v340[8:0], v4315[12:0]); // 3.0
    wire [17:0] v4316; shift_adder #(17, 15, 1, 1, 18, 3, 0) op_4316 (v1809[16:0], v1611[14:0], v4316[17:0]); // 3.0
    wire [13:0] v4317; shift_adder #(13, 13, 1, 1, 14, 0, 0) op_4317 (v2436[12:0], v813[12:0], v4317[13:0]); // 3.0
    wire [16:0] v4318; shift_adder #(13, 14, 1, 1, 17, 3, 0) op_4318 (v2437[12:0], v2438[13:0], v4318[16:0]); // 3.0
    wire [13:0] v4319; shift_adder #(12, 12, 1, 1, 14, 1, 0) op_4319 (v2341[11:0], v2072[11:0], v4319[13:0]); // 3.0
    wire [14:0] v4320; shift_adder #(13, 14, 1, 1, 15, 0, 0) op_4320 (v1670[12:0], v1790[13:0], v4320[14:0]); // 3.0
    wire [18:0] v4321; shift_adder #(18, 15, 1, 1, 19, 3, 0) op_4321 (v2439[17:0], v1880[14:0], v4321[18:0]); // 3.0
    wire [14:0] v4322; shift_adder #(12, 15, 1, 1, 15, 0, 0) op_4322 (v924[11:0], v2440[14:0], v4322[14:0]); // 3.0
    wire [14:0] v4323; shift_adder #(13, 12, 1, 1, 15, 2, 0) op_4323 (v2441[12:0], v1602[11:0], v4323[14:0]); // 3.0
    wire [14:0] v4324; shift_adder #(14, 12, 1, 1, 15, 2, 0) op_4324 (v1790[13:0], v825[11:0], v4324[14:0]); // 3.0
    wire [22:0] v4325; shift_adder #(14, 23, 1, 1, 23, -7, 0) op_4325 (v878[13:0], v1930[22:0], v4325[22:0]); // 3.0
    wire [13:0] v4326; shift_adder #(13, 10, 1, 1, 14, 2, 0) op_4326 (v2442[12:0], v2443[9:0], v4326[13:0]); // 3.0
    wire [20:0] v4327; shift_adder #(21, 13, 1, 1, 21, 6, 0) op_4327 (v1181[20:0], v2444[12:0], v4327[20:0]); // 3.0
    wire [20:0] v4328; shift_adder #(20, 11, 1, 1, 21, 8, 0) op_4328 (v2445[19:0], v772[10:0], v4328[20:0]); // 3.0
    wire [28:0] v4329; shift_adder #(28, 21, 1, 1, 29, 8, 0) op_4329 (v1022[27:0], v1596[20:0], v4329[28:0]); // 3.0
    wire [22:0] v4330; shift_adder #(11, 22, 1, 1, 23, -11, 0) op_4330 (v1581[10:0], v1664[21:0], v4330[22:0]); // 3.0
    wire [15:0] v4331; shift_adder #(13, 12, 1, 1, 16, 3, 0) op_4331 (v2446[12:0], v2447[11:0], v4331[15:0]); // 3.0
    wire [26:0] v4332; shift_adder #(25, 13, 1, 1, 27, 13, 0) op_4332 (v1935[24:0], v2390[12:0], v4332[26:0]); // 3.0
    wire [24:0] v4333; shift_adder #(18, 14, 1, 1, 25, -7, 0) op_4333 (v2289[17:0], v2412[13:0], v4333[24:0]); // 3.0
    wire [18:0] v4334; shift_adder #(19, 18, 1, 1, 19, 0, 0) op_4334 (v2448[18:0], v1835[17:0], v4334[18:0]); // 3.0
    wire [15:0] v4335; shift_adder #(11, 16, 1, 1, 16, -4, 0) op_4335 (v2234[10:0], v2449[15:0], v4335[15:0]); // 3.0
    wire [17:0] v4336; shift_adder #(15, 13, 1, 1, 18, 5, 0) op_4336 (v1084[14:0], v892[12:0], v4336[17:0]); // 3.0
    wire [20:0] v4337; shift_adder #(13, 19, 1, 1, 21, -7, 0) op_4337 (v2450[12:0], v1801[18:0], v4337[20:0]); // 3.0
    wire [24:0] v4338; shift_adder #(23, 25, 1, 1, 25, -1, 0) op_4338 (v1474[22:0], v1770[24:0], v4338[24:0]); // 3.0
    wire [23:0] v4339; shift_adder #(12, 23, 1, 1, 24, -11, 0) op_4339 (v1283[11:0], v2451[22:0], v4339[23:0]); // 3.0
    wire [15:0] v4340; shift_adder #(14, 15, 1, 1, 16, -1, 0) op_4340 (v2452[13:0], v2037[14:0], v4340[15:0]); // 3.0
    wire [19:0] v4341; shift_adder #(12, 19, 1, 1, 20, -6, 0) op_4341 (v2168[11:0], v2453[18:0], v4341[19:0]); // 3.0
    wire [36:0] v4342; shift_adder #(36, 18, 1, 1, 37, 19, 0) op_4342 (v2454[35:0], v1869[17:0], v4342[36:0]); // 3.0
    wire [19:0] v4343; shift_adder #(12, 19, 1, 1, 20, -7, 0) op_4343 (v2455[11:0], v1059[18:0], v4343[19:0]); // 3.0
    wire [13:0] v4344; shift_adder #(13, 12, 1, 1, 14, 1, 0) op_4344 (v1458[12:0], v1340[11:0], v4344[13:0]); // 3.0
    wire [17:0] v4345; shift_adder #(17, 15, 1, 1, 18, 3, 0) op_4345 (v1546[16:0], v2044[14:0], v4345[17:0]); // 3.0
    wire [12:0] v4346; shift_adder #(13, 12, 1, 1, 13, 0, 0) op_4346 (v2456[12:0], v1923[11:0], v4346[12:0]); // 3.0
    wire [21:0] v4347; shift_adder #(14, 21, 1, 1, 22, -7, 0) op_4347 (v2457[13:0], v998[20:0], v4347[21:0]); // 3.0
    wire [27:0] v4348; shift_adder #(17, 27, 1, 1, 28, -10, 0) op_4348 (v2458[16:0], v2359[26:0], v4348[27:0]); // 3.0
    wire [26:0] v4349; shift_adder #(26, 13, 1, 1, 27, 12, 0) op_4349 (v1881[25:0], v1872[12:0], v4349[26:0]); // 3.0
    wire [17:0] v4350; shift_adder #(15, 17, 1, 1, 18, -3, 1) op_4350 (v2022[14:0], v2173[16:0], v4350[17:0]); // 3.0
    wire [21:0] v4351; shift_adder #(21, 11, 1, 1, 22, 9, 0) op_4351 (v2206[20:0], v2459[10:0], v4351[21:0]); // 3.0
    wire [20:0] v4352; shift_adder #(13, 20, 1, 1, 21, -7, 0) op_4352 (v2010[12:0], v1384[19:0], v4352[20:0]); // 3.0
    wire [21:0] v4353; shift_adder #(22, 14, 1, 1, 22, 7, 0) op_4353 (v2460[21:0], v2461[13:0], v4353[21:0]); // 3.0
    wire [17:0] v4354; shift_adder #(15, 12, 1, 1, 18, 5, 0) op_4354 (v2243[14:0], v2108[11:0], v4354[17:0]); // 3.0
    wire [15:0] v4355; shift_adder #(16, 13, 1, 1, 16, 2, 0) op_4355 (v1557[15:0], v2462[12:0], v4355[15:0]); // 3.0
    wire [17:0] v4356; shift_adder #(17, 17, 1, 1, 18, -1, 0) op_4356 (v1023[16:0], v972[16:0], v4356[17:0]); // 3.0
    wire [17:0] v4357; shift_adder #(16, 17, 1, 1, 18, -1, 0) op_4357 (v1360[15:0], v2463[16:0], v4357[17:0]); // 3.0
    wire [14:0] v4358; shift_adder #(14, 13, 1, 1, 15, -1, 0) op_4358 (v2110[13:0], v2464[12:0], v4358[14:0]); // 3.0
    wire [13:0] v4359; shift_adder #(12, 13, 1, 1, 14, 0, 0) op_4359 (v1642[11:0], v1661[12:0], v4359[13:0]); // 3.0
    wire [13:0] v4360; shift_adder #(10, 14, 1, 1, 14, -2, 0) op_4360 (v2290[9:0], v1165[13:0], v4360[13:0]); // 3.0
    wire [16:0] v4361; shift_adder #(17, 14, 1, 1, 17, 1, 0) op_4361 (v2463[16:0], v1673[13:0], v4361[16:0]); // 3.0
    wire [18:0] v4362; shift_adder #(15, 18, 1, 1, 19, 1, 0) op_4362 (v1012[14:0], v2465[17:0], v4362[18:0]); // 3.0
    wire [14:0] v4363; shift_adder #(13, 13, 1, 1, 15, 1, 0) op_4363 (v2395[12:0], v1046[12:0], v4363[14:0]); // 3.0
    wire [16:0] v4364; shift_adder #(15, 14, 1, 1, 17, 2, 0) op_4364 (v2466[14:0], v1607[13:0], v4364[16:0]); // 3.0
    wire [13:0] v4365; shift_adder #(12, 12, 1, 1, 14, 1, 0) op_4365 (v1155[11:0], v1121[11:0], v4365[13:0]); // 3.0
    wire [22:0] v4366; shift_adder #(21, 11, 1, 1, 23, 12, 0) op_4366 (v943[20:0], v2467[10:0], v4366[22:0]); // 3.0
    wire [22:0] v4367; shift_adder #(11, 21, 1, 1, 23, -11, 0) op_4367 (v1523[10:0], v1403[20:0], v4367[22:0]); // 3.0
    wire [17:0] v4368; shift_adder #(17, 12, 1, 1, 18, 6, 0) op_4368 (v2468[16:0], v1082[11:0], v4368[17:0]); // 3.0
    wire [22:0] v4369; shift_adder #(22, 12, 1, 1, 23, 10, 0) op_4369 (v2460[21:0], v1031[11:0], v4369[22:0]); // 3.0
    wire [29:0] v4370; shift_adder #(12, 30, 1, 1, 30, -17, 0) op_4370 (v935[11:0], v2343[29:0], v4370[29:0]); // 3.0
    wire [14:0] v4371; shift_adder #(13, 12, 1, 1, 15, 2, 0) op_4371 (v1551[12:0], v1642[11:0], v4371[14:0]); // 3.0
    wire [27:0] v4372; shift_adder #(26, 19, 1, 1, 28, 9, 0) op_4372 (v1448[25:0], v2317[18:0], v4372[27:0]); // 3.0
    wire [22:0] v4373; shift_adder #(13, 22, 1, 1, 23, -8, 0) op_4373 (v2469[12:0], v844[21:0], v4373[22:0]); // 3.0
    wire [19:0] v4374; shift_adder #(11, 19, 1, 1, 20, -8, 0) op_4374 (v1517[10:0], v2470[18:0], v4374[19:0]); // 3.0
    wire [15:0] v4375; shift_adder #(12, 15, 1, 1, 16, -3, 0) op_4375 (v2471[11:0], v2117[14:0], v4375[15:0]); // 3.0
    wire [17:0] v4376; shift_adder #(18, 13, 1, 1, 18, 2, 0) op_4376 (v872[17:0], v1524[12:0], v4376[17:0]); // 3.0
    wire [12:0] v4377; shift_adder #(11, 12, 1, 1, 13, 0, 0) op_4377 (v2472[10:0], v2473[11:0], v4377[12:0]); // 3.0
    wire [20:0] v4378; shift_adder #(11, 21, 1, 1, 21, -7, 0) op_4378 (v1494[10:0], v2475[20:0], v4378[20:0]); // 3.0
    wire [26:0] v4379; shift_adder #(11, 26, 1, 1, 27, -15, 1) op_4379 (v251[10:0], v1838[25:0], v4379[26:0]); // 3.0
    wire [38:0] v4380; shift_adder #(33, 38, 1, 1, 39, -5, 0) op_4380 (v1779[32:0], v2476[37:0], v4380[38:0]); // 3.0
    wire [16:0] v4381; shift_adder #(16, 15, 1, 1, 17, 1, 0) op_4381 (v1929[15:0], v2414[14:0], v4381[16:0]); // 3.0
    wire [23:0] v4382; shift_adder #(16, 23, 1, 1, 24, -7, 0) op_4382 (v2150[15:0], v1842[22:0], v4382[23:0]); // 3.0
    wire [35:0] v4383; shift_adder #(34, 14, 1, 1, 36, -2, 1) op_4383 (v2477[33:0], v807[13:0], v4383[35:0]); // 3.0
    wire [36:0] v4384; shift_adder #(12, 12, 1, 1, 37, 25, 1) op_4384 (v2478[11:0], v438[11:0], v4384[36:0]); // 3.0
    wire [16:0] v4385; shift_adder #(13, 15, 1, 1, 17, -3, 0) op_4385 (v2375[12:0], v839[14:0], v4385[16:0]); // 3.0
    wire [12:0] v4386; shift_adder #(12, 12, 1, 1, 13, 1, 0) op_4386 (v1829[11:0], v929[11:0], v4386[12:0]); // 3.0
    wire [16:0] v4387; shift_adder #(15, 17, 1, 1, 17, 0, 0) op_4387 (v1535[14:0], v2479[16:0], v4387[16:0]); // 3.0
    wire [30:0] v4388; shift_adder #(29, 29, 1, 1, 31, -1, 0) op_4388 (v2153[28:0], v2480[28:0], v4388[30:0]); // 3.0
    wire [18:0] v4389; shift_adder #(18, 16, 1, 1, 19, 2, 0) op_4389 (v1150[17:0], v2271[15:0], v4389[18:0]); // 3.0
    wire [25:0] v4390; shift_adder #(26, 12, 1, 1, 26, 10, 0) op_4390 (v1791[25:0], v2481[11:0], v4390[25:0]); // 3.0
    wire [16:0] v4391; shift_adder #(15, 14, 1, 1, 17, 2, 0) op_4391 (v922[14:0], v2482[13:0], v4391[16:0]); // 3.0
    wire [16:0] v4392; shift_adder #(16, 11, 1, 1, 17, 4, 0) op_4392 (v2483[15:0], v1426[10:0], v4392[16:0]); // 3.0
    wire [24:0] v4393; shift_adder #(22, 25, 1, 1, 25, -2, 0) op_4393 (v1760[21:0], v1405[24:0], v4393[24:0]); // 3.0
    wire [19:0] v4394; shift_adder #(19, 17, 1, 1, 20, 2, 0) op_4394 (v1826[18:0], v2397[16:0], v4394[19:0]); // 3.0
    wire [20:0] v4395; shift_adder #(20, 20, 1, 1, 21, 0, 0) op_4395 (v2255[19:0], v1286[19:0], v4395[20:0]); // 3.0
    wire [24:0] v4396; shift_adder #(24, 19, 1, 1, 25, 5, 0) op_4396 (v2096[23:0], v2484[18:0], v4396[24:0]); // 3.0
    wire [16:0] v4397; shift_adder #(17, 10, 1, 1, 17, 5, 0) op_4397 (v2226[16:0], v2339[9:0], v4397[16:0]); // 3.0
    wire [20:0] v4398; shift_adder #(14, 20, 1, 1, 21, -5, 0) op_4398 (v1982[13:0], v2485[19:0], v4398[20:0]); // 3.0
    wire [19:0] v4399; shift_adder #(15, 18, 1, 1, 20, -4, 0) op_4399 (v1769[14:0], v1032[17:0], v4399[19:0]); // 3.0
    wire [13:0] v4400; shift_adder #(13, 13, 1, 1, 14, 0, 0) op_4400 (v2486[12:0], v2235[12:0], v4400[13:0]); // 3.0
    wire [14:0] v4401; shift_adder #(12, 13, 1, 1, 15, -2, 0) op_4401 (v1468[11:0], v2487[12:0], v4401[14:0]); // 3.0
    wire [22:0] v4402; shift_adder #(20, 23, 1, 1, 23, -1, 0) op_4402 (v2488[19:0], v1685[22:0], v4402[22:0]); // 3.0
    wire [26:0] v4403; shift_adder #(15, 27, 1, 1, 27, -9, 0) op_4403 (v1477[14:0], v2489[26:0], v4403[26:0]); // 3.0
    wire [23:0] v4404; shift_adder #(23, 15, 1, 1, 24, 8, 0) op_4404 (v1131[22:0], v2106[14:0], v4404[23:0]); // 3.0
    wire [26:0] v4405; shift_adder #(18, 26, 1, 1, 27, -8, 0) op_4405 (v2474[17:0], v2203[25:0], v4405[26:0]); // 3.0
    wire [27:0] v4406; shift_adder #(15, 27, 1, 1, 28, -13, 0) op_4406 (v1858[14:0], v2359[26:0], v4406[27:0]); // 3.0
    wire [22:0] v4407; shift_adder #(22, 14, 1, 1, 23, 9, 0) op_4407 (v1635[21:0], v2040[13:0], v4407[22:0]); // 3.0
    wire [19:0] v4408; shift_adder #(15, 19, 1, 1, 20, -2, 0) op_4408 (v1769[14:0], v2490[18:0], v4408[19:0]); // 3.0
    wire [17:0] v4409; shift_adder #(15, 17, 1, 1, 18, 1, 0) op_4409 (v2015[14:0], v1151[16:0], v4409[17:0]); // 3.0
    wire [17:0] v4410; shift_adder #(15, 12, 1, 1, 18, 5, 0) op_4410 (v1304[14:0], v2491[11:0], v4410[17:0]); // 3.0
    wire [14:0] v4411; shift_adder #(11, 14, 1, 1, 15, -2, 0) op_4411 (v2095[10:0], v2331[13:0], v4411[14:0]); // 3.0
    wire [21:0] v4412; shift_adder #(15, 22, 1, 1, 22, -6, 0) op_4412 (v2492[14:0], v1671[21:0], v4412[21:0]); // 3.0
    wire [28:0] v4413; shift_adder #(28, 17, 1, 1, 29, 11, 0) op_4413 (v2311[27:0], v2112[16:0], v4413[28:0]); // 3.0
    wire [21:0] v4414; shift_adder #(21, 19, 1, 1, 22, 2, 0) op_4414 (v1981[20:0], v2493[18:0], v4414[21:0]); // 3.0
    wire [27:0] v4415; shift_adder #(13, 27, 1, 1, 28, -14, 0) op_4415 (v1041[12:0], v933[26:0], v4415[27:0]); // 3.0
    wire [35:0] v4416; shift_adder #(13, 11, 1, 1, 36, 25, 1) op_4416 (v1660[12:0], v195[10:0], v4416[35:0]); // 3.0
    wire [23:0] v4417; shift_adder #(11, 24, 1, 1, 24, -12, 0) op_4417 (v2260[10:0], v1548[23:0], v4417[23:0]); // 3.0
    wire [15:0] v4418; shift_adder #(13, 16, 1, 1, 16, -2, 0) op_4418 (v2494[12:0], v2185[15:0], v4418[15:0]); // 3.0
    wire [14:0] v4419; shift_adder #(12, 12, 1, 1, 15, -3, 0) op_4419 (v2334[11:0], v2495[11:0], v4419[14:0]); // 3.0
    wire [12:0] v4420; shift_adder #(12, 12, 1, 1, 13, 0, 0) op_4420 (v1977[11:0], v1035[11:0], v4420[12:0]); // 3.0
    wire [16:0] v4421; shift_adder #(14, 17, 1, 1, 17, -2, 0) op_4421 (v2496[13:0], v1023[16:0], v4421[16:0]); // 3.0
    wire [17:0] v4422; shift_adder #(13, 17, 1, 1, 18, -4, 0) op_4422 (v2215[12:0], v2497[16:0], v4422[17:0]); // 3.0
    wire [14:0] v4423; shift_adder #(13, 13, 1, 1, 15, 2, 0) op_4423 (v1393[12:0], v2395[12:0], v4423[14:0]); // 3.0
    wire [14:0] v4424; shift_adder #(14, 15, 1, 1, 15, 0, 0) op_4424 (v1104[13:0], v2498[14:0], v4424[14:0]); // 3.0
    wire [13:0] v4425; shift_adder #(12, 13, 1, 1, 14, -1, 0) op_4425 (v2027[11:0], v2499[12:0], v4425[13:0]); // 3.0
    wire [16:0] v4426; shift_adder #(15, 13, 1, 1, 17, 4, 0) op_4426 (v2500[14:0], v1461[12:0], v4426[16:0]); // 3.0
    wire [17:0] v4427; shift_adder #(13, 17, 1, 1, 18, -4, 0) op_4427 (v2501[12:0], v1063[16:0], v4427[17:0]); // 3.0
    wire [18:0] v4428; shift_adder #(18, 18, 1, 1, 19, 1, 0) op_4428 (v2230[17:0], v1073[17:0], v4428[18:0]); // 3.0
    wire [34:0] v4429; shift_adder #(14, 35, 1, 1, 35, -20, 0) op_4429 (v2503[13:0], v2504[34:0], v4429[34:0]); // 3.0
    wire [19:0] v4430; shift_adder #(13, 19, 1, 1, 20, -6, 0) op_4430 (v1825[12:0], v1547[18:0], v4430[19:0]); // 3.0
    wire [33:0] v4431; shift_adder #(33, 11, 1, 1, 34, 21, 0) op_4431 (v2365[32:0], v2260[10:0], v4431[33:0]); // 3.0
    wire [30:0] v4432; shift_adder #(31, 17, 1, 1, 31, 12, 0) op_4432 (v2087[30:0], v952[16:0], v4432[30:0]); // 3.0
    wire [12:0] v4433; shift_adder #(13, 12, 1, 1, 13, 0, 0) op_4433 (v1336[12:0], v1376[11:0], v4433[12:0]); // 3.0
    wire [22:0] v4434; shift_adder #(17, 21, 1, 1, 23, -5, 0) op_4434 (v2505[16:0], v1926[20:0], v4434[22:0]); // 3.0
    wire [15:0] v4435; shift_adder #(12, 15, 1, 1, 16, -3, 0) op_4435 (v2506[11:0], v2060[14:0], v4435[15:0]); // 3.0
    wire [23:0] v4436; shift_adder #(15, 24, 1, 1, 24, -8, 0) op_4436 (v1767[14:0], v2041[23:0], v4436[23:0]); // 3.0
    wire [23:0] v4437; shift_adder #(23, 13, 1, 1, 24, 9, 0) op_4437 (v2507[22:0], v1781[12:0], v4437[23:0]); // 3.0
    wire [25:0] v4438; shift_adder #(26, 14, 1, 1, 26, 10, 0) op_4438 (v1042[25:0], v1538[13:0], v4438[25:0]); // 3.0
    wire [29:0] v4439; shift_adder #(29, 12, 1, 1, 30, 18, 0) op_4439 (v2508[28:0], v981[11:0], v4439[29:0]); // 3.0
    wire [12:0] v4440; shift_adder #(12, 12, 1, 1, 13, 1, 0) op_4440 (v794[11:0], v1443[11:0], v4440[12:0]); // 3.0
    wire [16:0] v4441; shift_adder #(14, 14, 1, 1, 17, -2, 0) op_4441 (v2509[13:0], v1939[13:0], v4441[16:0]); // 3.0
    wire [14:0] v4442; shift_adder #(12, 14, 1, 1, 15, -2, 0) op_4442 (v2135[11:0], v1165[13:0], v4442[14:0]); // 3.0
    wire [19:0] v4443; shift_adder #(14, 17, 1, 1, 20, -5, 0) op_4443 (v2510[13:0], v895[16:0], v4443[19:0]); // 3.0
    wire [15:0] v4444; shift_adder #(14, 13, 1, 1, 16, -2, 0) op_4444 (v2511[13:0], v2371[12:0], v4444[15:0]); // 3.0
    wire [20:0] v4445; shift_adder #(19, 16, 1, 1, 21, 5, 0) op_4445 (v2512[18:0], v2513[15:0], v4445[20:0]); // 4.0
    wire [24:0] v4446; shift_adder #(24, 22, 1, 1, 25, 1, 0) op_4446 (v2514[23:0], v2515[21:0], v4446[24:0]); // 4.0
    wire [22:0] v4447; shift_adder #(19, 22, 1, 1, 23, -3, 0) op_4447 (v2516[18:0], v2517[21:0], v4447[22:0]); // 4.0
    wire [24:0] v4448; shift_adder #(22, 24, 1, 1, 25, -2, 0) op_4448 (v2518[21:0], v2519[23:0], v4448[24:0]); // 4.0
    wire [25:0] v4449; shift_adder #(15, 26, 1, 1, 26, -8, 0) op_4449 (v781[14:0], v2520[25:0], v4449[25:0]); // 4.0
    wire [26:0] v4450; shift_adder #(25, 13, 1, 1, 27, 14, 0) op_4450 (v2521[24:0], v2522[12:0], v4450[26:0]); // 4.0
    wire [24:0] v4451; shift_adder #(15, 25, 1, 1, 25, -8, 0) op_4451 (v2523[14:0], v2524[24:0], v4451[24:0]); // 4.0
    wire [27:0] v4452; shift_adder #(13, 28, 1, 1, 28, -5, 1) op_4452 (v790[12:0], v2525[27:0], v4452[27:0]); // 4.0
    wire [24:0] v4453; shift_adder #(14, 24, 1, 1, 25, -10, 0) op_4453 (v2526[13:0], v2527[23:0], v4453[24:0]); // 4.0
    wire [17:0] v4454; shift_adder #(13, 17, 1, 1, 18, -5, 0) op_4454 (v2528[12:0], v2529[16:0], v4454[17:0]); // 4.0
    wire [27:0] v4455; shift_adder #(25, 23, 1, 1, 28, -3, 0) op_4455 (v796[24:0], v2530[22:0], v4455[27:0]); // 4.0
    wire [30:0] v4456; shift_adder #(28, 14, 1, 1, 31, 17, 0) op_4456 (v2531[27:0], v2532[13:0], v4456[30:0]); // 4.0
    wire [26:0] v4457; shift_adder #(8, 27, 1, 1, 27, -12, 0) op_4457 (v75[7:0], v2533[26:0], v4457[26:0]); // 4.0
    wire [16:0] v4458; shift_adder #(11, 14, 1, 1, 17, -6, 1) op_4458 (v191[10:0], v2534[13:0], v4458[16:0]); // 4.0
    wire [22:0] v4459; shift_adder #(22, 21, 1, 1, 23, 0, 0) op_4459 (v2535[21:0], v2536[20:0], v4459[22:0]); // 4.0
    wire [27:0] v4460; shift_adder #(13, 27, 1, 1, 28, -14, 0) op_4460 (v2537[12:0], v2538[26:0], v4460[27:0]); // 4.0
    wire [31:0] v4461; shift_adder #(31, 31, 1, 1, 32, 1, 0) op_4461 (v2539[30:0], v2540[30:0], v4461[31:0]); // 4.0
    wire [18:0] v4462; shift_adder #(17, 18, 1, 1, 19, 0, 0) op_4462 (v2541[16:0], v2542[17:0], v4462[18:0]); // 4.0
    wire [21:0] v4463; shift_adder #(18, 19, 1, 1, 22, -3, 0) op_4463 (v2543[17:0], v2544[18:0], v4463[21:0]); // 4.0
    wire [24:0] v4464; shift_adder #(8, 13, 1, 1, 25, 12, 0) op_4464 (v108[7:0], v2545[12:0], v4464[24:0]); // 4.0
    wire [14:0] v4465; shift_adder #(12, 15, 1, 1, 15, -2, 0) op_4465 (v2546[11:0], v2547[14:0], v4465[14:0]); // 4.0
    wire [15:0] v4466; shift_adder #(13, 15, 1, 1, 16, 0, 0) op_4466 (v2548[12:0], v2549[14:0], v4466[15:0]); // 4.0
    wire [27:0] v4467; shift_adder #(20, 27, 1, 1, 28, -8, 0) op_4467 (v2550[19:0], v2551[26:0], v4467[27:0]); // 4.0
    wire [23:0] v4468; shift_adder #(14, 24, 1, 1, 24, -9, 0) op_4468 (v2552[13:0], v2553[23:0], v4468[23:0]); // 4.0
    wire [19:0] v4469; shift_adder #(18, 15, 1, 1, 20, 5, 0) op_4469 (v2554[17:0], v2555[14:0], v4469[19:0]); // 4.0
    wire [26:0] v4470; shift_adder #(10, 18, 1, 1, 27, -17, 0) op_4470 (v235[9:0], v2556[17:0], v4470[26:0]); // 4.0
    wire [28:0] v4471; shift_adder #(17, 28, 1, 1, 29, -11, 0) op_4471 (v2557[16:0], v2558[27:0], v4471[28:0]); // 4.0
    wire [20:0] v4472; shift_adder #(17, 20, 1, 1, 21, -2, 0) op_4472 (v2559[16:0], v2560[19:0], v4472[20:0]); // 4.0
    wire [22:0] v4473; shift_adder #(17, 23, 1, 1, 23, -4, 0) op_4473 (v2561[16:0], v2562[22:0], v4473[22:0]); // 4.0
    wire [21:0] v4474; shift_adder #(8, 22, 1, 1, 22, 0, 1) op_4474 (v78[7:0], v2563[21:0], v4474[21:0]); // 4.0
    wire [17:0] v4475; shift_adder #(16, 18, 1, 1, 18, 0, 0) op_4475 (v2564[15:0], v2565[17:0], v4475[17:0]); // 4.0
    wire [30:0] v4476; shift_adder #(16, 31, 1, 1, 31, -13, 0) op_4476 (v2566[15:0], v2567[30:0], v4476[30:0]); // 4.0
    wire [28:0] v4477; shift_adder #(29, 18, 1, 1, 29, 10, 0) op_4477 (v2568[28:0], v2569[17:0], v4477[28:0]); // 4.0
    wire [34:0] v4478; shift_adder #(18, 34, 1, 1, 35, -15, 0) op_4478 (v2570[17:0], v2571[33:0], v4478[34:0]); // 4.0
    wire [16:0] v4479; shift_adder #(13, 16, 1, 1, 17, -3, 0) op_4479 (v2572[12:0], v2573[15:0], v4479[16:0]); // 4.0
    wire [14:0] v4480; shift_adder #(14, 13, 1, 1, 15, 0, 0) op_4480 (v2574[13:0], v2575[12:0], v4480[14:0]); // 4.0
    wire [31:0] v4481; shift_adder #(31, 19, 1, 1, 32, 12, 0) op_4481 (v2576[30:0], v2577[18:0], v4481[31:0]); // 4.0
    wire [22:0] v4482; shift_adder #(15, 22, 1, 1, 23, 1, 1) op_4482 (v2578[14:0], v868[21:0], v4482[22:0]); // 4.0
    wire [19:0] v4483; shift_adder #(17, 18, 1, 1, 20, -2, 0) op_4483 (v2579[16:0], v2580[17:0], v4483[19:0]); // 4.0
    wire [18:0] v4484; shift_adder #(14, 18, 1, 1, 19, -5, 0) op_4484 (v249[13:0], v2581[17:0], v4484[18:0]); // 4.0
    wire [18:0] v4485; shift_adder #(18, 15, 1, 1, 19, 0, 0) op_4485 (v2582[17:0], v2583[14:0], v4485[18:0]); // 4.0
    wire [18:0] v4486; shift_adder #(12, 19, 1, 1, 19, -6, 0) op_4486 (v879[11:0], v2584[18:0], v4486[18:0]); // 4.0
    wire [21:0] v4487; shift_adder #(19, 14, 1, 1, 22, 7, 0) op_4487 (v2585[18:0], v2586[13:0], v4487[21:0]); // 4.0
    wire [24:0] v4488; shift_adder #(14, 22, 1, 1, 25, 3, 0) op_4488 (v290[13:0], v2587[21:0], v4488[24:0]); // 4.0
    wire [20:0] v4489; shift_adder #(13, 18, 1, 1, 21, -7, 0) op_4489 (v2588[12:0], v2589[17:0], v4489[20:0]); // 4.0
    wire [21:0] v4490; shift_adder #(20, 17, 1, 1, 22, 4, 0) op_4490 (v2590[19:0], v2591[16:0], v4490[21:0]); // 4.0
    wire [21:0] v4491; shift_adder #(8, 21, 1, 1, 22, 1, 0) op_4491 (v104[7:0], v2592[20:0], v4491[21:0]); // 4.0
    wire [15:0] v4492; shift_adder #(11, 15, 1, 1, 16, -5, 0) op_4492 (v215[10:0], v2593[14:0], v4492[15:0]); // 4.0
    wire [16:0] v4493; shift_adder #(15, 16, 1, 1, 17, -1, 0) op_4493 (v2594[14:0], v2595[15:0], v4493[16:0]); // 4.0
    wire [19:0] v4494; shift_adder #(8, 20, 1, 1, 20, -3, 0) op_4494 (v97[7:0], v2596[19:0], v4494[19:0]); // 4.0
    wire [19:0] v4495; shift_adder #(18, 15, 1, 1, 20, 5, 0) op_4495 (v2597[17:0], v2598[14:0], v4495[19:0]); // 4.0
    wire [19:0] v4496; shift_adder #(18, 17, 1, 1, 20, 3, 0) op_4496 (v2599[17:0], v2600[16:0], v4496[19:0]); // 4.0
    wire [20:0] v4497; shift_adder #(20, 20, 1, 1, 21, 1, 0) op_4497 (v2601[19:0], v2602[19:0], v4497[20:0]); // 4.0
    wire [26:0] v4498; shift_adder #(27, 22, 1, 1, 27, 2, 0) op_4498 (v2603[26:0], v2604[21:0], v4498[26:0]); // 4.0
    wire [22:0] v4499; shift_adder #(22, 20, 1, 1, 23, 2, 0) op_4499 (v2605[21:0], v2606[19:0], v4499[22:0]); // 4.0
    wire [28:0] v4500; shift_adder #(28, 17, 1, 1, 29, 11, 0) op_4500 (v2607[27:0], v2608[16:0], v4500[28:0]); // 4.0
    wire [34:0] v4501; shift_adder #(13, 35, 1, 1, 35, -3, 1) op_4501 (v149[12:0], v2609[34:0], v4501[34:0]); // 4.0
    wire [22:0] v4502; shift_adder #(22, 18, 1, 1, 23, 3, 0) op_4502 (v2610[21:0], v2611[17:0], v4502[22:0]); // 4.0
    wire [19:0] v4503; shift_adder #(13, 18, 1, 1, 20, -6, 0) op_4503 (v2612[12:0], v2613[17:0], v4503[19:0]); // 4.0
    wire [16:0] v4504; shift_adder #(15, 16, 1, 1, 17, 1, 0) op_4504 (v318[14:0], v2614[15:0], v4504[16:0]); // 4.0
    wire [22:0] v4505; shift_adder #(17, 23, 1, 1, 23, -3, 0) op_4505 (v2615[16:0], v2616[22:0], v4505[22:0]); // 4.0
    wire [25:0] v4506; shift_adder #(8, 25, 1, 1, 26, -17, 0) op_4506 (v65[7:0], v2617[24:0], v4506[25:0]); // 4.0
    wire [19:0] v4507; shift_adder #(19, 15, 1, 1, 20, 4, 0) op_4507 (v2618[18:0], v2619[14:0], v4507[19:0]); // 4.0
    wire [26:0] v4508; shift_adder #(27, 22, 1, 1, 27, 2, 0) op_4508 (v2620[26:0], v2621[21:0], v4508[26:0]); // 4.0
    wire [19:0] v4509; shift_adder #(11, 15, 1, 1, 20, 5, 0) op_4509 (v229[10:0], v2622[14:0], v4509[19:0]); // 4.0
    wire [27:0] v4510; shift_adder #(27, 26, 1, 1, 28, 1, 0) op_4510 (v2623[26:0], v2624[25:0], v4510[27:0]); // 4.0
    wire [30:0] v4511; shift_adder #(11, 15, 1, 1, 31, -20, 0) op_4511 (v245[10:0], v2625[14:0], v4511[30:0]); // 4.0
    wire [19:0] v4512; shift_adder #(18, 19, 1, 1, 20, 0, 0) op_4512 (v2626[17:0], v2627[18:0], v4512[19:0]); // 4.0
    wire [22:0] v4513; shift_adder #(21, 22, 1, 1, 23, -1, 0) op_4513 (v2628[20:0], v2629[21:0], v4513[22:0]); // 4.0
    wire [33:0] v4514; shift_adder #(21, 34, 1, 1, 34, -12, 0) op_4514 (v2630[20:0], v2631[33:0], v4514[33:0]); // 4.0
    wire [27:0] v4515; shift_adder #(26, 18, 1, 1, 28, 9, 0) op_4515 (v2632[25:0], v2633[17:0], v4515[27:0]); // 4.0
    wire [25:0] v4516; shift_adder #(8, 26, 1, 1, 26, -1, 0) op_4516 (v82[7:0], v2634[25:0], v4516[25:0]); // 4.0
    wire [35:0] v4517; shift_adder #(18, 35, 1, 1, 36, -16, 0) op_4517 (v2635[17:0], v2636[34:0], v4517[35:0]); // 4.0
    wire [16:0] v4518; shift_adder #(16, 14, 1, 1, 17, -1, 0) op_4518 (v2637[15:0], v2638[13:0], v4518[16:0]); // 4.0
    wire [17:0] v4519; shift_adder #(16, 18, 1, 1, 18, -1, 0) op_4519 (v2639[15:0], v2640[17:0], v4519[17:0]); // 4.0
    wire [17:0] v4520; shift_adder #(17, 17, 1, 1, 18, 0, 0) op_4520 (v2641[16:0], v2642[16:0], v4520[17:0]); // 4.0
    wire [18:0] v4521; shift_adder #(17, 18, 1, 1, 19, -2, 0) op_4521 (v2643[16:0], v2644[17:0], v4521[18:0]); // 4.0
    wire [21:0] v4522; shift_adder #(18, 21, 1, 1, 22, -3, 0) op_4522 (v2645[17:0], v2646[20:0], v4522[21:0]); // 4.0
    wire [20:0] v4523; shift_adder #(20, 21, 1, 1, 21, 0, 0) op_4523 (v2647[19:0], v2648[20:0], v4523[20:0]); // 4.0
    wire [18:0] v4524; shift_adder #(16, 18, 1, 1, 19, -2, 0) op_4524 (v2649[15:0], v2650[17:0], v4524[18:0]); // 4.0
    wire [15:0] v4525; shift_adder #(14, 15, 1, 1, 16, 0, 0) op_4525 (v2651[13:0], v2652[14:0], v4525[15:0]); // 4.0
    wire [19:0] v4526; shift_adder #(8, 19, 1, 1, 20, 1, 0) op_4526 (v120[7:0], v2653[18:0], v4526[19:0]); // 4.0
    wire [28:0] v4527; shift_adder #(19, 28, 1, 1, 29, -9, 0) op_4527 (v2654[18:0], v2655[27:0], v4527[28:0]); // 4.0
    wire [26:0] v4528; shift_adder #(18, 26, 1, 1, 27, -8, 0) op_4528 (v2656[17:0], v2624[25:0], v4528[26:0]); // 4.0
    wire [19:0] v4529; shift_adder #(17, 19, 1, 1, 20, -2, 0) op_4529 (v2657[16:0], v2658[18:0], v4529[19:0]); // 4.0
    wire [38:0] v4530; shift_adder #(38, 31, 1, 1, 39, 7, 0) op_4530 (v2659[37:0], v2660[30:0], v4530[38:0]); // 4.0
    wire [37:0] v4531; shift_adder #(16, 26, 1, 1, 38, 12, 1) op_4531 (v2661[15:0], v988[25:0], v4531[37:0]); // 4.0
    wire [27:0] v4532; shift_adder #(27, 19, 1, 1, 28, 9, 0) op_4532 (v2551[26:0], v2662[18:0], v4532[27:0]); // 4.0
    wire [14:0] v4533; shift_adder #(14, 14, 1, 1, 15, -1, 0) op_4533 (v2663[13:0], v2664[13:0], v4533[14:0]); // 4.0
    wire [23:0] v4534; shift_adder #(16, 23, 1, 1, 24, -6, 0) op_4534 (v2665[15:0], v2666[22:0], v4534[23:0]); // 4.0
    wire [22:0] v4535; shift_adder #(23, 19, 1, 1, 23, 2, 0) op_4535 (v2667[22:0], v2668[18:0], v4535[22:0]); // 4.0
    wire [23:0] v4536; shift_adder #(23, 19, 1, 1, 24, 3, 0) op_4536 (v2669[22:0], v2670[18:0], v4536[23:0]); // 4.0
    wire [22:0] v4537; shift_adder #(11, 19, 1, 1, 23, 4, 0) op_4537 (v199[10:0], v2671[18:0], v4537[22:0]); // 4.0
    wire [24:0] v4538; shift_adder #(14, 23, 1, 1, 25, -10, 0) op_4538 (v2672[13:0], v2673[22:0], v4538[24:0]); // 4.0
    wire [13:0] v4539; shift_adder #(10, 13, 1, 1, 14, 1, 1) op_4539 (v366[9:0], v2674[12:0], v4539[13:0]); // 4.0
    wire [24:0] v4540; shift_adder #(8, 25, 1, 1, 25, -3, 1) op_4540 (v126[7:0], v2675[24:0], v4540[24:0]); // 4.0
    wire [22:0] v4541; shift_adder #(17, 23, 1, 1, 23, -5, 0) op_4541 (v2676[16:0], v2677[22:0], v4541[22:0]); // 4.0
    wire [25:0] v4542; shift_adder #(19, 26, 1, 1, 26, -4, 0) op_4542 (v2678[18:0], v2679[25:0], v4542[25:0]); // 4.0
    wire [29:0] v4543; shift_adder #(16, 30, 1, 1, 30, -12, 0) op_4543 (v2680[15:0], v2681[29:0], v4543[29:0]); // 4.0
    wire [26:0] v4544; shift_adder #(8, 22, 1, 1, 27, 5, 1) op_4544 (v65[7:0], v2682[21:0], v4544[26:0]); // 4.0
    wire [22:0] v4545; shift_adder #(11, 23, 1, 1, 23, -11, 0) op_4545 (v377[10:0], v2683[22:0], v4545[22:0]); // 4.0
    wire [25:0] v4546; shift_adder #(25, 16, 1, 1, 26, 8, 0) op_4546 (v2684[24:0], v2685[15:0], v4546[25:0]); // 4.0
    wire [16:0] v4547; shift_adder #(8, 17, 1, 1, 17, -5, 1) op_4547 (v100[7:0], v2686[16:0], v4547[16:0]); // 4.0
    wire [34:0] v4548; shift_adder #(31, 34, 1, 1, 35, -3, 1) op_4548 (v381[30:0], v2687[33:0], v4548[34:0]); // 4.0
    wire [30:0] v4549; shift_adder #(31, 14, 1, 1, 31, 15, 0) op_4549 (v2688[30:0], v2689[13:0], v4549[30:0]); // 4.0
    wire [19:0] v4550; shift_adder #(18, 18, 1, 1, 20, 1, 0) op_4550 (v2690[17:0], v2691[17:0], v4550[19:0]); // 4.0
    wire [26:0] v4551; shift_adder #(11, 14, 1, 1, 27, 13, 0) op_4551 (v334[10:0], v2692[13:0], v4551[26:0]); // 4.0
    wire [22:0] v4552; shift_adder #(8, 22, 1, 1, 23, -13, 1) op_4552 (v71[7:0], v2693[21:0], v4552[22:0]); // 4.0
    wire [20:0] v4553; shift_adder #(15, 20, 1, 1, 21, -4, 0) op_4553 (v2694[14:0], v2695[19:0], v4553[20:0]); // 4.0
    wire [19:0] v4554; shift_adder #(17, 19, 1, 1, 20, -2, 0) op_4554 (v2696[16:0], v2697[18:0], v4554[19:0]); // 4.0
    wire [22:0] v4555; shift_adder #(22, 21, 1, 1, 23, 0, 0) op_4555 (v2698[21:0], v2699[20:0], v4555[22:0]); // 4.0
    wire [31:0] v4556; shift_adder #(8, 26, 1, 1, 32, 6, 0) op_4556 (v80[7:0], v2700[25:0], v4556[31:0]); // 4.0
    wire [27:0] v4557; shift_adder #(26, 25, 1, 1, 28, -2, 0) op_4557 (v2701[25:0], v2702[24:0], v4557[27:0]); // 4.0
    wire [16:0] v4558; shift_adder #(14, 15, 1, 1, 17, -3, 0) op_4558 (v2703[13:0], v2704[14:0], v4558[16:0]); // 4.0
    wire [38:0] v4559; shift_adder #(15, 13, 1, 1, 39, 26, 1) op_4559 (v2705[14:0], v1048[12:0], v4559[38:0]); // 4.0
    wire [34:0] v4560; shift_adder #(26, 34, 1, 1, 35, -8, 0) op_4560 (v2706[25:0], v2707[33:0], v4560[34:0]); // 4.0
    wire [16:0] v4561; shift_adder #(16, 15, 1, 1, 17, 1, 0) op_4561 (v2708[15:0], v2709[14:0], v4561[16:0]); // 4.0
    wire [16:0] v4562; shift_adder #(15, 16, 1, 1, 17, -2, 0) op_4562 (v2710[14:0], v2711[15:0], v4562[16:0]); // 4.0
    wire [31:0] v4563; shift_adder #(12, 32, 1, 1, 32, -7, 1) op_4563 (v304[11:0], v2712[31:0], v4563[31:0]); // 4.0
    wire [33:0] v4564; shift_adder #(25, 33, 1, 1, 34, -8, 0) op_4564 (v2702[24:0], v2713[32:0], v4564[33:0]); // 4.0
    wire [25:0] v4565; shift_adder #(23, 25, 1, 1, 26, -2, 0) op_4565 (v2714[22:0], v2715[24:0], v4565[25:0]); // 4.0
    wire [36:0] v4566; shift_adder #(21, 36, 1, 1, 37, -14, 0) op_4566 (v2716[20:0], v2717[35:0], v4566[36:0]); // 4.0
    wire [22:0] v4567; shift_adder #(23, 14, 1, 1, 23, 7, 0) op_4567 (v2718[22:0], v2719[13:0], v4567[22:0]); // 4.0
    wire [16:0] v4568; shift_adder #(16, 15, 1, 1, 17, -1, 0) op_4568 (v2720[15:0], v2721[14:0], v4568[16:0]); // 4.0
    wire [20:0] v4569; shift_adder #(19, 20, 1, 1, 21, -1, 0) op_4569 (v2722[18:0], v2723[19:0], v4569[20:0]); // 4.0
    wire [27:0] v4570; shift_adder #(21, 27, 1, 1, 28, -7, 0) op_4570 (v2630[20:0], v2724[26:0], v4570[27:0]); // 4.0
    wire [18:0] v4571; shift_adder #(13, 18, 1, 1, 19, -5, 0) op_4571 (v2725[12:0], v2726[17:0], v4571[18:0]); // 4.0
    wire [18:0] v4572; shift_adder #(18, 13, 1, 1, 19, 6, 0) op_4572 (v2727[17:0], v2728[12:0], v4572[18:0]); // 4.0
    wire [18:0] v4573; shift_adder #(14, 16, 1, 1, 19, -4, 0) op_4573 (v2729[13:0], v2730[15:0], v4573[18:0]); // 4.0
    wire [15:0] v4574; shift_adder #(15, 14, 1, 1, 16, 0, 0) op_4574 (v2731[14:0], v2732[13:0], v4574[15:0]); // 4.0
    wire [26:0] v4575; shift_adder #(12, 27, 1, 1, 27, -13, 0) op_4575 (v2733[11:0], v2734[26:0], v4575[26:0]); // 4.0
    wire [21:0] v4576; shift_adder #(8, 21, 1, 1, 22, -12, 0) op_4576 (v105[7:0], v2735[20:0], v4576[21:0]); // 4.0
    wire [28:0] v4577; shift_adder #(27, 21, 1, 1, 29, 8, 0) op_4577 (v2736[26:0], v2737[20:0], v4577[28:0]); // 4.0
    wire [30:0] v4578; shift_adder #(30, 18, 1, 1, 31, 13, 0) op_4578 (v2738[29:0], v2726[17:0], v4578[30:0]); // 4.0
    wire [26:0] v4579; shift_adder #(20, 25, 1, 1, 27, -6, 0) op_4579 (v2739[19:0], v2740[24:0], v4579[26:0]); // 4.0
    wire [32:0] v4580; shift_adder #(31, 32, 1, 1, 33, 1, 0) op_4580 (v2741[30:0], v2742[31:0], v4580[32:0]); // 4.0
    wire [28:0] v4581; shift_adder #(28, 18, 1, 1, 29, 10, 0) op_4581 (v2743[27:0], v2744[17:0], v4581[28:0]); // 4.0
    wire [21:0] v4582; shift_adder #(13, 21, 1, 1, 22, -6, 0) op_4582 (v2745[12:0], v2746[20:0], v4582[21:0]); // 4.0
    wire [16:0] v4583; shift_adder #(15, 14, 1, 1, 17, 2, 0) op_4583 (v2747[14:0], v2748[13:0], v4583[16:0]); // 4.0
    wire [19:0] v4584; shift_adder #(18, 15, 1, 1, 20, 5, 0) op_4584 (v2749[17:0], v2750[14:0], v4584[19:0]); // 4.0
    wire [21:0] v4585; shift_adder #(21, 18, 1, 1, 22, 3, 0) op_4585 (v2751[20:0], v2752[17:0], v4585[21:0]); // 4.0
    wire [36:0] v4586; shift_adder #(16, 35, 1, 1, 37, -21, 0) op_4586 (v2753[15:0], v2754[34:0], v4586[36:0]); // 4.0
    wire [26:0] v4587; shift_adder #(20, 26, 1, 1, 27, -7, 0) op_4587 (v2755[19:0], v2756[25:0], v4587[26:0]); // 4.0
    wire [16:0] v4588; shift_adder #(15, 15, 1, 1, 17, -1, 0) op_4588 (v2757[14:0], v2758[14:0], v4588[16:0]); // 4.0
    wire [19:0] v4589; shift_adder #(20, 16, 1, 1, 20, 1, 0) op_4589 (v2759[19:0], v2760[15:0], v4589[19:0]); // 4.0
    wire [18:0] v4590; shift_adder #(18, 14, 1, 1, 19, 3, 0) op_4590 (v2761[17:0], v2762[13:0], v4590[18:0]); // 4.0
    wire [17:0] v4591; shift_adder #(15, 18, 1, 1, 18, -2, 0) op_4591 (v2763[14:0], v2764[17:0], v4591[17:0]); // 4.0
    wire [17:0] v4592; shift_adder #(15, 17, 1, 1, 18, 1, 0) op_4592 (v2765[14:0], v2766[16:0], v4592[17:0]); // 4.0
    wire [20:0] v4593; shift_adder #(21, 17, 1, 1, 21, 3, 0) op_4593 (v2767[20:0], v2768[16:0], v4593[20:0]); // 4.0
    wire [22:0] v4594; shift_adder #(19, 22, 1, 1, 23, -4, 0) op_4594 (v2769[18:0], v2770[21:0], v4594[22:0]); // 4.0
    wire [24:0] v4595; shift_adder #(23, 24, 1, 1, 25, -1, 0) op_4595 (v2771[22:0], v2772[23:0], v4595[24:0]); // 4.0
    wire [32:0] v4596; shift_adder #(11, 19, 1, 1, 33, 14, 1) op_4596 (v329[10:0], v2773[18:0], v4596[32:0]); // 4.0
    wire [19:0] v4597; shift_adder #(19, 14, 1, 1, 20, 6, 0) op_4597 (v2774[18:0], v2775[13:0], v4597[19:0]); // 4.0
    wire [30:0] v4598; shift_adder #(14, 31, 1, 1, 31, -14, 0) op_4598 (v2776[13:0], v2777[30:0], v4598[30:0]); // 4.0
    wire [25:0] v4599; shift_adder #(24, 21, 1, 1, 26, 5, 0) op_4599 (v2778[23:0], v2779[20:0], v4599[25:0]); // 4.0
    wire [24:0] v4600; shift_adder #(24, 24, 1, 1, 25, -1, 0) op_4600 (v2780[23:0], v2781[23:0], v4600[24:0]); // 4.0
    wire [30:0] v4601; shift_adder #(18, 31, 1, 1, 31, -12, 0) op_4601 (v2599[17:0], v2782[30:0], v4601[30:0]); // 4.0
    wire [24:0] v4602; shift_adder #(17, 14, 1, 1, 25, 11, 0) op_4602 (v1146[16:0], v2783[13:0], v4602[24:0]); // 4.0
    wire [26:0] v4603; shift_adder #(25, 24, 1, 1, 27, 2, 0) op_4603 (v2784[24:0], v2785[23:0], v4603[26:0]); // 4.0
    wire [19:0] v4604; shift_adder #(15, 19, 1, 1, 20, -4, 0) op_4604 (v922[14:0], v2786[18:0], v4604[19:0]); // 4.0
    wire [16:0] v4605; shift_adder #(16, 14, 1, 1, 17, 2, 0) op_4605 (v2787[15:0], v2788[13:0], v4605[16:0]); // 4.0
    wire [29:0] v4606; shift_adder #(28, 17, 1, 1, 30, 12, 0) op_4606 (v2789[27:0], v2790[16:0], v4606[29:0]); // 4.0
    wire [37:0] v4607; shift_adder #(19, 37, 1, 1, 38, -19, 0) op_4607 (v2791[18:0], v2792[36:0], v4607[37:0]); // 4.0
    wire [16:0] v4608; shift_adder #(14, 15, 1, 1, 17, -2, 0) op_4608 (v2793[13:0], v2794[14:0], v4608[16:0]); // 4.0
    wire [17:0] v4609; shift_adder #(15, 15, 1, 1, 18, -3, 0) op_4609 (v2795[14:0], v2796[14:0], v4609[17:0]); // 4.0
    wire [18:0] v4610; shift_adder #(8, 19, 1, 1, 19, -6, 0) op_4610 (v111[7:0], v2797[18:0], v4610[18:0]); // 4.0
    wire [28:0] v4611; shift_adder #(29, 26, 1, 1, 29, 0, 0) op_4611 (v2798[28:0], v2799[25:0], v4611[28:0]); // 4.0
    wire [31:0] v4612; shift_adder #(32, 17, 1, 1, 32, 12, 0) op_4612 (v2800[31:0], v2801[16:0], v4612[31:0]); // 4.0
    wire [28:0] v4613; shift_adder #(11, 19, 1, 1, 29, 10, 1) op_4613 (v195[10:0], v2802[18:0], v4613[28:0]); // 4.0
    wire [25:0] v4614; shift_adder #(25, 17, 1, 1, 26, 7, 0) op_4614 (v2803[24:0], v2804[16:0], v4614[25:0]); // 4.0
    wire [17:0] v4615; shift_adder #(18, 14, 1, 1, 18, 2, 0) op_4615 (v2805[17:0], v2806[13:0], v4615[17:0]); // 4.0
    wire [21:0] v4616; shift_adder #(22, 17, 1, 1, 22, 1, 0) op_4616 (v2807[21:0], v2643[16:0], v4616[21:0]); // 4.0
    wire [21:0] v4617; shift_adder #(22, 18, 1, 1, 22, 3, 0) op_4617 (v2808[21:0], v2809[17:0], v4617[21:0]); // 4.0
    wire [16:0] v4618; shift_adder #(14, 16, 1, 1, 17, -3, 0) op_4618 (v2810[13:0], v2811[15:0], v4618[16:0]); // 4.0
    wire [32:0] v4619; shift_adder #(32, 24, 1, 1, 33, 8, 0) op_4619 (v2812[31:0], v2813[23:0], v4619[32:0]); // 4.0
    wire [35:0] v4620; shift_adder #(35, 24, 1, 1, 36, 11, 0) op_4620 (v2814[34:0], v2815[23:0], v4620[35:0]); // 4.0
    wire [35:0] v4621; shift_adder #(35, 14, 1, 1, 36, 22, 0) op_4621 (v2816[34:0], v2817[13:0], v4621[35:0]); // 4.0
    wire [32:0] v4622; shift_adder #(14, 32, 1, 1, 33, -18, 0) op_4622 (v2818[13:0], v2819[31:0], v4622[32:0]); // 4.0
    wire [17:0] v4623; shift_adder #(11, 18, 1, 1, 18, 0, 1) op_4623 (v821[10:0], v2820[17:0], v4623[17:0]); // 4.0
    wire [29:0] v4624; shift_adder #(28, 22, 1, 1, 30, 8, 0) op_4624 (v2821[27:0], v2822[21:0], v4624[29:0]); // 4.0
    wire [30:0] v4625; shift_adder #(27, 29, 1, 1, 31, -3, 0) op_4625 (v2823[26:0], v2824[28:0], v4625[30:0]); // 4.0
    wire [30:0] v4626; shift_adder #(31, 12, 1, 1, 31, 5, 1) op_4626 (v2825[30:0], v1199[11:0], v4626[30:0]); // 4.0
    wire [25:0] v4627; shift_adder #(23, 25, 1, 1, 26, -2, 0) op_4627 (v2826[22:0], v2827[24:0], v4627[25:0]); // 4.0
    wire [22:0] v4628; shift_adder #(23, 14, 1, 1, 23, 7, 0) op_4628 (v2828[22:0], v2829[13:0], v4628[22:0]); // 4.0
    wire [20:0] v4629; shift_adder #(15, 20, 1, 1, 21, -4, 0) op_4629 (v2795[14:0], v2830[19:0], v4629[20:0]); // 4.0
    wire [24:0] v4630; shift_adder #(16, 22, 1, 1, 25, -8, 0) op_4630 (v2831[15:0], v2832[21:0], v4630[24:0]); // 4.0
    wire [29:0] v4631; shift_adder #(8, 30, 1, 1, 30, -1, 1) op_4631 (v90[7:0], v2833[29:0], v4631[29:0]); // 4.0
    wire [19:0] v4632; shift_adder #(20, 18, 1, 1, 20, 1, 0) op_4632 (v2834[19:0], v2835[17:0], v4632[19:0]); // 4.0
    wire [19:0] v4633; shift_adder #(13, 20, 1, 1, 20, -5, 0) op_4633 (v2836[12:0], v2837[19:0], v4633[19:0]); // 4.0
    wire [23:0] v4634; shift_adder #(22, 17, 1, 1, 24, 7, 0) op_4634 (v2838[21:0], v2676[16:0], v4634[23:0]); // 4.0
    wire [27:0] v4635; shift_adder #(15, 26, 1, 1, 28, -12, 0) op_4635 (v2839[14:0], v2840[25:0], v4635[27:0]); // 4.0
    wire [29:0] v4636; shift_adder #(21, 29, 1, 1, 30, -7, 0) op_4636 (v2841[20:0], v2842[28:0], v4636[29:0]); // 4.0
    wire [21:0] v4637; shift_adder #(8, 22, 1, 1, 22, -3, 0) op_4637 (v78[7:0], v2843[21:0], v4637[21:0]); // 4.0
    wire [31:0] v4638; shift_adder #(30, 21, 1, 1, 32, 10, 0) op_4638 (v2844[29:0], v2845[20:0], v4638[31:0]); // 4.0
    wire [22:0] v4639; shift_adder #(21, 19, 1, 1, 23, 3, 0) op_4639 (v2846[20:0], v2847[18:0], v4639[22:0]); // 4.0
    wire [14:0] v4640; shift_adder #(14, 14, 1, 1, 15, 0, 0) op_4640 (v2848[13:0], v2849[13:0], v4640[14:0]); // 4.0
    wire [18:0] v4641; shift_adder #(15, 18, 1, 1, 19, -2, 0) op_4641 (v2850[14:0], v2851[17:0], v4641[18:0]); // 4.0
    wire [28:0] v4642; shift_adder #(9, 22, 1, 1, 29, -19, 1) op_4642 (v231[8:0], v2852[21:0], v4642[28:0]); // 4.0
    wire [30:0] v4643; shift_adder #(30, 25, 1, 1, 31, 5, 0) op_4643 (v2853[29:0], v2854[24:0], v4643[30:0]); // 4.0
    wire [25:0] v4644; shift_adder #(21, 24, 1, 1, 26, -4, 0) op_4644 (v2855[20:0], v2778[23:0], v4644[25:0]); // 4.0
    wire [23:0] v4645; shift_adder #(8, 24, 1, 1, 24, -6, 0) op_4645 (v67[7:0], v2856[23:0], v4645[23:0]); // 4.0
    wire [30:0] v4646; shift_adder #(13, 25, 1, 1, 31, -18, 0) op_4646 (v1097[12:0], v2857[24:0], v4646[30:0]); // 4.0
    wire [31:0] v4647; shift_adder #(31, 20, 1, 1, 32, 12, 0) op_4647 (v2858[30:0], v2602[19:0], v4647[31:0]); // 4.0
    wire [16:0] v4648; shift_adder #(16, 13, 1, 1, 17, 2, 0) op_4648 (v2859[15:0], v2860[12:0], v4648[16:0]); // 4.0
    wire [32:0] v4649; shift_adder #(8, 22, 1, 1, 33, 11, 0) op_4649 (v113[7:0], v2862[21:0], v4649[32:0]); // 4.0
    wire [18:0] v4650; shift_adder #(15, 16, 1, 1, 19, 2, 0) op_4650 (v471[14:0], v2863[15:0], v4650[18:0]); // 4.0
    wire [29:0] v4651; shift_adder #(29, 15, 1, 1, 30, 14, 0) op_4651 (v2864[28:0], v2865[14:0], v4651[29:0]); // 4.0
    wire [25:0] v4652; shift_adder #(12, 19, 1, 1, 26, -14, 1) op_4652 (v1178[11:0], v2866[18:0], v4652[25:0]); // 4.0
    wire [33:0] v4653; shift_adder #(32, 28, 1, 1, 34, 5, 0) op_4653 (v2867[31:0], v2868[27:0], v4653[33:0]); // 4.0
    wire [18:0] v4654; shift_adder #(18, 13, 1, 1, 19, 5, 0) op_4654 (v2569[17:0], v2869[12:0], v4654[18:0]); // 4.0
    wire [16:0] v4655; shift_adder #(17, 13, 1, 1, 17, 3, 0) op_4655 (v2870[16:0], v2869[12:0], v4655[16:0]); // 4.0
    wire [18:0] v4656; shift_adder #(14, 18, 1, 1, 19, -4, 0) op_4656 (v2871[13:0], v2872[17:0], v4656[18:0]); // 4.0
    wire [34:0] v4657; shift_adder #(20, 34, 1, 1, 35, -14, 0) op_4657 (v2873[19:0], v2874[33:0], v4657[34:0]); // 4.0
    wire [16:0] v4658; shift_adder #(17, 13, 1, 1, 17, 2, 0) op_4658 (v2875[16:0], v2876[12:0], v4658[16:0]); // 4.0
    wire [39:0] v4659; shift_adder #(16, 17, 1, 1, 40, -24, 1) op_4659 (v2877[15:0], v2878[16:0], v4659[39:0]); // 4.0
    wire [28:0] v4660; shift_adder #(13, 28, 1, 1, 29, -15, 0) op_4660 (v2879[12:0], v2880[27:0], v4660[28:0]); // 4.0
    wire [25:0] v4661; shift_adder #(24, 13, 1, 1, 26, 12, 0) op_4661 (v2881[23:0], v2537[12:0], v4661[25:0]); // 4.0
    wire [27:0] v4662; shift_adder #(8, 28, 1, 1, 28, -10, 0) op_4662 (v88[7:0], v2882[27:0], v4662[27:0]); // 4.0
    wire [30:0] v4663; shift_adder #(8, 29, 1, 1, 31, -22, 1) op_4663 (v91[7:0], v2883[28:0], v4663[30:0]); // 4.0
    wire [23:0] v4664; shift_adder #(22, 17, 1, 1, 24, 7, 0) op_4664 (v2698[21:0], v2884[16:0], v4664[23:0]); // 4.0
    wire [21:0] v4665; shift_adder #(21, 19, 1, 1, 22, 1, 0) op_4665 (v2885[20:0], v2585[18:0], v4665[21:0]); // 4.0
    wire [28:0] v4666; shift_adder #(24, 27, 1, 1, 29, -4, 0) op_4666 (v2886[23:0], v2887[26:0], v4666[28:0]); // 4.0
    wire [31:0] v4667; shift_adder #(27, 31, 1, 1, 32, -3, 0) op_4667 (v2888[26:0], v2889[30:0], v4667[31:0]); // 4.0
    wire [29:0] v4668; shift_adder #(29, 17, 1, 1, 30, 11, 0) op_4668 (v2890[28:0], v2891[16:0], v4668[29:0]); // 4.0
    wire [15:0] v4669; shift_adder #(13, 15, 1, 1, 16, -2, 0) op_4669 (v2892[12:0], v2893[14:0], v4669[15:0]); // 4.0
    wire [16:0] v4670; shift_adder #(15, 16, 1, 1, 17, -2, 0) op_4670 (v2894[14:0], v2895[15:0], v4670[16:0]); // 4.0
    wire [23:0] v4671; shift_adder #(11, 17, 1, 1, 24, -13, 0) op_4671 (v323[10:0], v2768[16:0], v4671[23:0]); // 4.0
    wire [20:0] v4672; shift_adder #(13, 21, 1, 1, 21, -7, 0) op_4672 (v2896[12:0], v2897[20:0], v4672[20:0]); // 4.0
    wire [24:0] v4673; shift_adder #(25, 24, 1, 1, 25, 0, 0) op_4673 (v2898[24:0], v2899[23:0], v4673[24:0]); // 4.0
    wire [22:0] v4674; shift_adder #(22, 22, 1, 1, 23, 0, 0) op_4674 (v2832[21:0], v2900[21:0], v4674[22:0]); // 4.0
    wire [21:0] v4675; shift_adder #(14, 21, 1, 1, 22, -7, 0) op_4675 (v2901[13:0], v2902[20:0], v4675[21:0]); // 4.0
    wire [17:0] v4676; shift_adder #(14, 17, 1, 1, 18, -4, 0) op_4676 (v2903[13:0], v2904[16:0], v4676[17:0]); // 4.0
    wire [25:0] v4677; shift_adder #(24, 16, 1, 1, 26, 9, 0) op_4677 (v2905[23:0], v2906[15:0], v4677[25:0]); // 4.0
    wire [15:0] v4678; shift_adder #(14, 14, 1, 1, 16, 2, 0) op_4678 (v2907[13:0], v2908[13:0], v4678[15:0]); // 4.0
    wire [20:0] v4679; shift_adder #(18, 21, 1, 1, 21, -2, 0) op_4679 (v2726[17:0], v2909[20:0], v4679[20:0]); // 4.0
    wire [20:0] v4680; shift_adder #(16, 18, 1, 1, 21, 3, 0) op_4680 (v2910[15:0], v2911[17:0], v4680[20:0]); // 4.0
    wire [22:0] v4681; shift_adder #(15, 23, 1, 1, 23, -5, 0) op_4681 (v2912[14:0], v2913[22:0], v4681[22:0]); // 4.0
    wire [23:0] v4682; shift_adder #(15, 23, 1, 1, 24, -7, 0) op_4682 (v2914[14:0], v2915[22:0], v4682[23:0]); // 4.0
    wire [19:0] v4683; shift_adder #(16, 18, 1, 1, 20, -3, 0) op_4683 (v2916[15:0], v2917[17:0], v4683[19:0]); // 4.0
    wire [19:0] v4684; shift_adder #(16, 18, 1, 1, 20, -3, 0) op_4684 (v2918[15:0], v2919[17:0], v4684[19:0]); // 4.0
    wire [19:0] v4685; shift_adder #(17, 19, 1, 1, 20, -2, 0) op_4685 (v2920[16:0], v2774[18:0], v4685[19:0]); // 4.0
    wire [18:0] v4686; shift_adder #(18, 17, 1, 1, 19, 1, 0) op_4686 (v2921[17:0], v2922[16:0], v4686[18:0]); // 4.0
    wire [32:0] v4687; shift_adder #(33, 22, 1, 1, 33, 8, 0) op_4687 (v2923[32:0], v2924[21:0], v4687[32:0]); // 4.0
    wire [28:0] v4688; shift_adder #(8, 26, 1, 1, 29, -20, 1) op_4688 (v82[7:0], v2925[25:0], v4688[28:0]); // 4.0
    wire [28:0] v4689; shift_adder #(28, 21, 1, 1, 29, 7, 0) op_4689 (v2926[27:0], v2927[20:0], v4689[28:0]); // 4.0
    wire [33:0] v4690; shift_adder #(8, 33, 1, 1, 34, -24, 0) op_4690 (v72[7:0], v2928[32:0], v4690[33:0]); // 4.0
    wire [32:0] v4691; shift_adder #(13, 33, 1, 1, 33, -18, 0) op_4691 (v2929[12:0], v2930[32:0], v4691[32:0]); // 4.0
    wire [23:0] v4692; shift_adder #(24, 17, 1, 1, 24, 6, 0) op_4692 (v2931[23:0], v2932[16:0], v4692[23:0]); // 4.0
    wire [19:0] v4693; shift_adder #(17, 19, 1, 1, 20, -2, 0) op_4693 (v2657[16:0], v2933[18:0], v4693[19:0]); // 4.0
    wire [15:0] v4694; shift_adder #(15, 15, 1, 1, 16, 0, 0) op_4694 (v2934[14:0], v2935[14:0], v4694[15:0]); // 4.0
    wire [16:0] v4695; shift_adder #(11, 14, 1, 1, 17, 3, 1) op_4695 (v154[10:0], v2664[13:0], v4695[16:0]); // 4.0
    wire [33:0] v4696; shift_adder #(34, 25, 1, 1, 34, 8, 0) op_4696 (v2936[33:0], v2937[24:0], v4696[33:0]); // 4.0
    wire [16:0] v4697; shift_adder #(16, 13, 1, 1, 17, 3, 0) op_4697 (v2938[15:0], v2939[12:0], v4697[16:0]); // 4.0
    wire [23:0] v4698; shift_adder #(22, 20, 1, 1, 24, 3, 0) op_4698 (v2940[21:0], v2647[19:0], v4698[23:0]); // 4.0
    wire [34:0] v4699; shift_adder #(25, 35, 1, 1, 35, -9, 0) op_4699 (v2941[24:0], v2942[34:0], v4699[34:0]); // 4.0
    wire [26:0] v4700; shift_adder #(26, 13, 1, 1, 27, 13, 0) op_4700 (v2943[25:0], v2944[12:0], v4700[26:0]); // 4.0
    wire [24:0] v4701; shift_adder #(25, 23, 1, 1, 25, 0, 0) op_4701 (v2945[24:0], v2530[22:0], v4701[24:0]); // 4.0
    wire [29:0] v4702; shift_adder #(29, 23, 1, 1, 30, 6, 0) op_4702 (v2946[28:0], v2947[22:0], v4702[29:0]); // 4.0
    wire [20:0] v4703; shift_adder #(19, 16, 1, 1, 21, 5, 0) op_4703 (v2948[18:0], v2949[15:0], v4703[20:0]); // 4.0
    wire [23:0] v4704; shift_adder #(23, 20, 1, 1, 24, 3, 0) op_4704 (v2950[22:0], v2951[19:0], v4704[23:0]); // 4.0
    wire [23:0] v4705; shift_adder #(12, 16, 1, 1, 24, 8, 1) op_4705 (v457[11:0], v2952[15:0], v4705[23:0]); // 4.0
    wire [14:0] v4706; shift_adder #(14, 13, 1, 1, 15, 1, 0) op_4706 (v2953[13:0], v2954[12:0], v4706[14:0]); // 4.0
    wire [20:0] v4707; shift_adder #(21, 13, 1, 1, 21, 6, 0) op_4707 (v2955[20:0], v2956[12:0], v4707[20:0]); // 4.0
    wire [17:0] v4708; shift_adder #(17, 15, 1, 1, 18, 0, 0) op_4708 (v2957[16:0], v2958[14:0], v4708[17:0]); // 4.0
    wire [30:0] v4709; shift_adder #(25, 31, 1, 1, 31, -4, 0) op_4709 (v2959[24:0], v2960[30:0], v4709[30:0]); // 4.0
    wire [14:0] v4710; shift_adder #(8, 14, 1, 1, 15, -5, 1) op_4710 (v115[7:0], v2961[13:0], v4710[14:0]); // 4.0
    wire [18:0] v4711; shift_adder #(11, 15, 1, 1, 19, -8, 1) op_4711 (v299[10:0], v2893[14:0], v4711[18:0]); // 4.0
    wire [25:0] v4712; shift_adder #(25, 21, 1, 1, 26, 3, 0) op_4712 (v2962[24:0], v2646[20:0], v4712[25:0]); // 4.0
    wire [29:0] v4713; shift_adder #(15, 30, 1, 1, 30, -13, 0) op_4713 (v2963[14:0], v2964[29:0], v4713[29:0]); // 4.0
    wire [31:0] v4714; shift_adder #(11, 13, 1, 1, 32, -21, 1) op_4714 (v237[10:0], v2965[12:0], v4714[31:0]); // 4.0
    wire [16:0] v4715; shift_adder #(16, 15, 1, 1, 17, 1, 0) op_4715 (v2966[15:0], v2967[14:0], v4715[16:0]); // 4.0
    wire [38:0] v4716; shift_adder #(38, 16, 1, 1, 39, 22, 0) op_4716 (v2969[37:0], v2970[15:0], v4716[38:0]); // 4.0
    wire [40:0] v4717; shift_adder #(31, 18, 1, 1, 41, -10, 1) op_4717 (v2971[30:0], v2972[17:0], v4717[40:0]); // 4.0
    wire [18:0] v4718; shift_adder #(12, 17, 1, 1, 19, -7, 0) op_4718 (v2973[11:0], v2974[16:0], v4718[18:0]); // 4.0
    wire [14:0] v4719; shift_adder #(8, 13, 1, 1, 15, 2, 0) op_4719 (v76[7:0], v2975[12:0], v4719[14:0]); // 4.0
    wire [16:0] v4720; shift_adder #(15, 16, 1, 1, 17, -1, 0) op_4720 (v2976[14:0], v2977[15:0], v4720[16:0]); // 4.0
    wire [16:0] v4721; shift_adder #(8, 14, 1, 1, 17, 3, 0) op_4721 (v91[7:0], v2978[13:0], v4721[16:0]); // 4.0
    wire [16:0] v4722; shift_adder #(15, 16, 1, 1, 17, 0, 0) op_4722 (v2979[14:0], v2980[15:0], v4722[16:0]); // 4.0
    wire [22:0] v4723; shift_adder #(20, 15, 1, 1, 23, 7, 0) op_4723 (v2981[19:0], v2982[14:0], v4723[22:0]); // 4.0
    wire [19:0] v4724; shift_adder #(14, 20, 1, 1, 20, 0, 1) op_4724 (v2983[13:0], v515[19:0], v4724[19:0]); // 4.0
    wire [15:0] v4725; shift_adder #(14, 15, 1, 1, 16, 0, 0) op_4725 (v2762[13:0], v2984[14:0], v4725[15:0]); // 4.0
    wire [21:0] v4726; shift_adder #(17, 14, 1, 1, 22, -5, 1) op_4726 (v972[16:0], v2985[13:0], v4726[21:0]); // 4.0
    wire [17:0] v4727; shift_adder #(17, 15, 1, 1, 18, 2, 0) op_4727 (v2986[16:0], v2987[14:0], v4727[17:0]); // 4.0
    wire [25:0] v4728; shift_adder #(23, 26, 1, 1, 26, 0, 0) op_4728 (v2988[22:0], v2989[25:0], v4728[25:0]); // 4.0
    wire [19:0] v4729; shift_adder #(19, 17, 1, 1, 20, 2, 0) op_4729 (v2990[18:0], v2615[16:0], v4729[19:0]); // 4.0
    wire [16:0] v4730; shift_adder #(14, 16, 1, 1, 17, -2, 0) op_4730 (v2991[13:0], v2992[15:0], v4730[16:0]); // 4.0
    wire [25:0] v4731; shift_adder #(22, 25, 1, 1, 26, -3, 0) op_4731 (v2993[21:0], v2994[24:0], v4731[25:0]); // 4.0
    wire [21:0] v4732; shift_adder #(8, 22, 1, 1, 22, -5, 0) op_4732 (v90[7:0], v2995[21:0], v4732[21:0]); // 4.0
    wire [22:0] v4733; shift_adder #(15, 22, 1, 1, 23, -6, 0) op_4733 (v2996[14:0], v2997[21:0], v4733[22:0]); // 4.0
    wire [23:0] v4734; shift_adder #(21, 19, 1, 1, 24, 5, 0) op_4734 (v2998[20:0], v2999[18:0], v4734[23:0]); // 4.0
    wire [22:0] v4735; shift_adder #(16, 22, 1, 1, 23, -6, 0) op_4735 (v3000[15:0], v3001[21:0], v4735[22:0]); // 4.0
    wire [30:0] v4736; shift_adder #(14, 31, 1, 1, 31, -16, 0) op_4736 (v3002[13:0], v3003[30:0], v4736[30:0]); // 4.0
    wire [27:0] v4737; shift_adder #(26, 26, 1, 1, 28, -2, 0) op_4737 (v3004[25:0], v3005[25:0], v4737[27:0]); // 4.0
    wire [22:0] v4738; shift_adder #(17, 22, 1, 1, 23, -4, 0) op_4738 (v3006[16:0], v3007[21:0], v4738[22:0]); // 4.0
    wire [35:0] v4739; shift_adder #(35, 24, 1, 1, 36, 11, 0) op_4739 (v3008[34:0], v3009[23:0], v4739[35:0]); // 4.0
    wire [22:0] v4740; shift_adder #(17, 20, 1, 1, 23, -6, 0) op_4740 (v3010[16:0], v3011[19:0], v4740[22:0]); // 4.0
    wire [17:0] v4741; shift_adder #(17, 14, 1, 1, 18, 3, 0) op_4741 (v3012[16:0], v3013[13:0], v4741[17:0]); // 4.0
    wire [23:0] v4742; shift_adder #(11, 24, 1, 1, 24, -10, 0) op_4742 (v176[10:0], v3014[23:0], v4742[23:0]); // 4.0
    wire [16:0] v4743; shift_adder #(13, 15, 1, 1, 17, -3, 0) op_4743 (v3015[12:0], v3016[14:0], v4743[16:0]); // 4.0
    wire [18:0] v4744; shift_adder #(18, 18, 1, 1, 19, 0, 0) op_4744 (v3017[17:0], v3018[17:0], v4744[18:0]); // 4.0
    wire [15:0] v4745; shift_adder #(8, 16, 1, 1, 16, 0, 0) op_4745 (v118[7:0], v3019[15:0], v4745[15:0]); // 4.0
    wire [25:0] v4746; shift_adder #(26, 20, 1, 1, 26, 4, 0) op_4746 (v3020[25:0], v3021[19:0], v4746[25:0]); // 4.0
    wire [34:0] v4747; shift_adder #(34, 20, 1, 1, 35, 13, 0) op_4747 (v3022[33:0], v3023[19:0], v4747[34:0]); // 4.0
    wire [33:0] v4748; shift_adder #(13, 26, 1, 1, 34, 8, 1) op_4748 (v3024[12:0], v1428[25:0], v4748[33:0]); // 4.0
    wire [26:0] v4749; shift_adder #(11, 16, 1, 1, 27, 11, 0) op_4749 (v197[10:0], v3025[15:0], v4749[26:0]); // 4.0
    wire [34:0] v4750; shift_adder #(33, 14, 1, 1, 35, 20, 0) op_4750 (v3026[32:0], v3027[13:0], v4750[34:0]); // 4.0
    wire [38:0] v4751; shift_adder #(14, 38, 1, 1, 39, -23, 0) op_4751 (v3028[13:0], v3029[37:0], v4751[38:0]); // 4.0
    wire [37:0] v4752; shift_adder #(14, 15, 1, 1, 38, -24, 1) op_4752 (v3030[13:0], v3031[14:0], v4752[37:0]); // 4.0
    wire [34:0] v4753; shift_adder #(15, 34, 1, 1, 35, -19, 0) op_4753 (v3032[14:0], v3033[33:0], v4753[34:0]); // 4.0
    wire [31:0] v4754; shift_adder #(31, 26, 1, 1, 32, 4, 0) op_4754 (v3034[30:0], v3035[25:0], v4754[31:0]); // 4.0
    wire [22:0] v4755; shift_adder #(22, 22, 1, 1, 23, 0, 0) op_4755 (v3036[21:0], v3037[21:0], v4755[22:0]); // 4.0
    wire [28:0] v4756; shift_adder #(16, 27, 1, 1, 29, -12, 0) op_4756 (v3038[15:0], v3039[26:0], v4756[28:0]); // 4.0
    wire [24:0] v4757; shift_adder #(24, 15, 1, 1, 25, 9, 0) op_4757 (v3040[23:0], v2555[14:0], v4757[24:0]); // 4.0
    wire [27:0] v4758; shift_adder #(27, 18, 1, 1, 28, 9, 0) op_4758 (v3041[26:0], v3042[17:0], v4758[27:0]); // 4.0
    wire [28:0] v4759; shift_adder #(26, 27, 1, 1, 29, -3, 0) op_4759 (v3043[25:0], v3044[26:0], v4759[28:0]); // 4.0
    wire [24:0] v4760; shift_adder #(15, 23, 1, 1, 25, -9, 0) op_4760 (v3045[14:0], v3046[22:0], v4760[24:0]); // 4.0
    wire [22:0] v4761; shift_adder #(11, 21, 1, 1, 23, 2, 1) op_4761 (v169[10:0], v3047[20:0], v4761[22:0]); // 4.0
    wire [23:0] v4762; shift_adder #(24, 14, 1, 1, 24, 9, 0) op_4762 (v3048[23:0], v3049[13:0], v4762[23:0]); // 4.0
    wire [24:0] v4763; shift_adder #(11, 22, 1, 1, 25, -14, 0) op_4763 (v323[10:0], v3050[21:0], v4763[24:0]); // 4.0
    wire [25:0] v4764; shift_adder #(21, 24, 1, 1, 26, -5, 0) op_4764 (v3051[20:0], v3052[23:0], v4764[25:0]); // 4.0
    wire [20:0] v4765; shift_adder #(13, 17, 1, 1, 21, -7, 0) op_4765 (v3053[12:0], v3054[16:0], v4765[20:0]); // 4.0
    wire [20:0] v4766; shift_adder #(13, 20, 1, 1, 21, -6, 0) op_4766 (v2572[12:0], v3055[19:0], v4766[20:0]); // 4.0
    wire [24:0] v4767; shift_adder #(17, 24, 1, 1, 25, -6, 0) op_4767 (v3056[16:0], v3057[23:0], v4767[24:0]); // 4.0
    wire [20:0] v4768; shift_adder #(16, 20, 1, 1, 21, -4, 0) op_4768 (v3058[15:0], v3059[19:0], v4768[20:0]); // 4.0
    wire [23:0] v4769; shift_adder #(24, 14, 1, 1, 24, 9, 0) op_4769 (v3060[23:0], v3061[13:0], v4769[23:0]); // 4.0
    wire [24:0] v4770; shift_adder #(23, 22, 1, 1, 25, 2, 0) op_4770 (v3062[22:0], v3063[21:0], v4770[24:0]); // 4.0
    wire [28:0] v4771; shift_adder #(27, 17, 1, 1, 29, 11, 0) op_4771 (v3064[26:0], v3065[16:0], v4771[28:0]); // 4.0
    wire [20:0] v4772; shift_adder #(20, 18, 1, 1, 21, 2, 0) op_4772 (v3066[19:0], v3067[17:0], v4772[20:0]); // 4.0
    wire [20:0] v4773; shift_adder #(18, 20, 1, 1, 21, 0, 0) op_4773 (v3068[17:0], v3069[19:0], v4773[20:0]); // 4.0
    wire [29:0] v4774; shift_adder #(28, 22, 1, 1, 30, 8, 0) op_4774 (v3070[27:0], v2563[21:0], v4774[29:0]); // 4.0
    wire [32:0] v4775; shift_adder #(32, 22, 1, 1, 33, 9, 0) op_4775 (v3071[31:0], v3072[21:0], v4775[32:0]); // 4.0
    wire [25:0] v4776; shift_adder #(26, 18, 1, 1, 26, 6, 0) op_4776 (v3073[25:0], v3074[17:0], v4776[25:0]); // 4.0
    wire [32:0] v4777; shift_adder #(27, 32, 1, 1, 33, -6, 0) op_4777 (v3075[26:0], v3076[31:0], v4777[32:0]); // 4.0
    wire [32:0] v4778; shift_adder #(27, 32, 1, 1, 33, -4, 0) op_4778 (v3077[26:0], v3078[31:0], v4778[32:0]); // 4.0
    wire [24:0] v4779; shift_adder #(17, 24, 1, 1, 25, -7, 0) op_4779 (v2804[16:0], v3079[23:0], v4779[24:0]); // 4.0
    wire [38:0] v4780; shift_adder #(36, 38, 1, 1, 39, -1, 0) op_4780 (v3080[35:0], v3081[37:0], v4780[38:0]); // 4.0
    wire [14:0] v4781; shift_adder #(13, 13, 1, 1, 15, 1, 0) op_4781 (v3082[12:0], v3083[12:0], v4781[14:0]); // 4.0
    wire [16:0] v4782; shift_adder #(13, 15, 1, 1, 17, 2, 0) op_4782 (v3084[12:0], v3085[14:0], v4782[16:0]); // 4.0
    wire [17:0] v4783; shift_adder #(15, 16, 1, 1, 18, -2, 0) op_4783 (v3086[14:0], v3087[15:0], v4783[17:0]); // 4.0
    wire [19:0] v4784; shift_adder #(14, 19, 1, 1, 20, -5, 0) op_4784 (v3088[13:0], v3089[18:0], v4784[19:0]); // 4.0
    wire [29:0] v4785; shift_adder #(29, 16, 1, 1, 30, 13, 0) op_4785 (v3090[28:0], v3091[15:0], v4785[29:0]); // 4.0
    wire [22:0] v4786; shift_adder #(21, 19, 1, 1, 23, 3, 0) op_4786 (v3092[20:0], v2847[18:0], v4786[22:0]); // 4.0
    wire [18:0] v4787; shift_adder #(13, 19, 1, 1, 19, -3, 0) op_4787 (v3093[12:0], v3094[18:0], v4787[18:0]); // 4.0
    wire [15:0] v4788; shift_adder #(15, 14, 1, 1, 16, -1, 0) op_4788 (v3095[14:0], v3096[13:0], v4788[15:0]); // 4.0
    wire [17:0] v4789; shift_adder #(10, 17, 1, 1, 18, 1, 0) op_4789 (v549[9:0], v2920[16:0], v4789[17:0]); // 4.0
    wire [19:0] v4790; shift_adder #(18, 19, 1, 1, 20, -1, 0) op_4790 (v3097[17:0], v3098[18:0], v4790[19:0]); // 4.0
    wire [25:0] v4791; shift_adder #(26, 12, 1, 1, 26, 12, 0) op_4791 (v3099[25:0], v3100[11:0], v4791[25:0]); // 4.0
    wire [17:0] v4792; shift_adder #(15, 15, 1, 1, 18, -3, 0) op_4792 (v3101[14:0], v3102[14:0], v4792[17:0]); // 4.0
    wire [23:0] v4793; shift_adder #(20, 24, 1, 1, 24, -3, 0) op_4793 (v3103[19:0], v3104[23:0], v4793[23:0]); // 4.0
    wire [16:0] v4794; shift_adder #(12, 15, 1, 1, 17, 2, 1) op_4794 (v1462[11:0], v3105[14:0], v4794[16:0]); // 4.0
    wire [14:0] v4795; shift_adder #(14, 13, 1, 1, 15, 1, 0) op_4795 (v3106[13:0], v3107[12:0], v4795[14:0]); // 4.0
    wire [21:0] v4796; shift_adder #(22, 18, 1, 1, 22, 3, 0) op_4796 (v2518[21:0], v3108[17:0], v4796[21:0]); // 4.0
    wire [22:0] v4797; shift_adder #(21, 22, 1, 1, 23, -1, 0) op_4797 (v3109[20:0], v3110[21:0], v4797[22:0]); // 4.0
    wire [16:0] v4798; shift_adder #(16, 16, 1, 1, 17, -1, 0) op_4798 (v3111[15:0], v3112[15:0], v4798[16:0]); // 4.0
    wire [25:0] v4799; shift_adder #(18, 25, 1, 1, 26, -7, 0) op_4799 (v2851[17:0], v2827[24:0], v4799[25:0]); // 4.0
    wire [28:0] v4800; shift_adder #(12, 21, 1, 1, 29, -17, 1) op_4800 (v552[11:0], v3113[20:0], v4800[28:0]); // 4.0
    wire [24:0] v4801; shift_adder #(15, 24, 1, 1, 25, -9, 0) op_4801 (v3114[14:0], v3115[23:0], v4801[24:0]); // 4.0
    wire [28:0] v4802; shift_adder #(29, 19, 1, 1, 29, 9, 0) op_4802 (v3116[28:0], v3117[18:0], v4802[28:0]); // 4.0
    wire [28:0] v4803; shift_adder #(28, 13, 1, 1, 29, 14, 0) op_4803 (v3118[27:0], v3119[12:0], v4803[28:0]); // 4.0
    wire [26:0] v4804; shift_adder #(26, 24, 1, 1, 27, -1, 0) op_4804 (v3120[25:0], v3121[23:0], v4804[26:0]); // 4.0
    wire [24:0] v4805; shift_adder #(15, 23, 1, 1, 25, -10, 0) op_4805 (v3122[14:0], v3123[22:0], v4805[24:0]); // 4.0
    wire [21:0] v4806; shift_adder #(16, 12, 1, 1, 22, -6, 0) op_4806 (v3124[15:0], v1261[11:0], v4806[21:0]); // 4.0
    wire [23:0] v4807; shift_adder #(12, 17, 1, 1, 24, 7, 0) op_4807 (v552[11:0], v3125[16:0], v4807[23:0]); // 4.0
    wire [28:0] v4808; shift_adder #(22, 28, 1, 1, 29, -5, 0) op_4808 (v3126[21:0], v3127[27:0], v4808[28:0]); // 4.0
    wire [19:0] v4809; shift_adder #(15, 18, 1, 1, 20, -5, 0) op_4809 (v3045[14:0], v3128[17:0], v4809[19:0]); // 4.0
    wire [19:0] v4810; shift_adder #(18, 18, 1, 1, 20, 1, 0) op_4810 (v3129[17:0], v3130[17:0], v4810[19:0]); // 4.0
    wire [19:0] v4811; shift_adder #(18, 18, 1, 1, 20, 2, 0) op_4811 (v2820[17:0], v3131[17:0], v4811[19:0]); // 4.0
    wire [25:0] v4812; shift_adder #(21, 25, 1, 1, 26, -3, 0) op_4812 (v3132[20:0], v3133[24:0], v4812[25:0]); // 4.0
    wire [25:0] v4813; shift_adder #(25, 14, 1, 1, 26, 12, 0) op_4813 (v3134[24:0], v3135[13:0], v4813[25:0]); // 4.0
    wire [20:0] v4814; shift_adder #(14, 20, 1, 1, 21, -5, 0) op_4814 (v3136[13:0], v3137[19:0], v4814[20:0]); // 4.0
    wire [27:0] v4815; shift_adder #(8, 23, 1, 1, 28, -19, 0) op_4815 (v66[7:0], v3138[22:0], v4815[27:0]); // 4.0
    wire [24:0] v4816; shift_adder #(24, 14, 1, 1, 25, 10, 0) op_4816 (v3139[23:0], v3140[13:0], v4816[24:0]); // 4.0
    wire [18:0] v4817; shift_adder #(19, 17, 1, 1, 19, 0, 0) op_4817 (v3141[18:0], v3142[16:0], v4817[18:0]); // 4.0
    wire [22:0] v4818; shift_adder #(19, 21, 1, 1, 23, -3, 0) op_4818 (v3143[18:0], v3144[20:0], v4818[22:0]); // 4.0
    wire [23:0] v4819; shift_adder #(8, 19, 1, 1, 24, 5, 0) op_4819 (v98[7:0], v3145[18:0], v4819[23:0]); // 4.0
    wire [22:0] v4820; shift_adder #(15, 21, 1, 1, 23, -8, 0) op_4820 (v3146[14:0], v3147[20:0], v4820[22:0]); // 4.0
    wire [19:0] v4821; shift_adder #(20, 14, 1, 1, 20, 4, 0) op_4821 (v3103[19:0], v3148[13:0], v4821[19:0]); // 4.0
    wire [24:0] v4822; shift_adder #(14, 25, 1, 1, 25, -10, 0) op_4822 (v3149[13:0], v3150[24:0], v4822[24:0]); // 4.0
    wire [18:0] v4823; shift_adder #(13, 17, 1, 1, 19, -5, 0) op_4823 (v3151[12:0], v3152[16:0], v4823[18:0]); // 4.0
    wire [21:0] v4824; shift_adder #(22, 19, 1, 1, 22, 0, 0) op_4824 (v3153[21:0], v3154[18:0], v4824[21:0]); // 4.0
    wire [18:0] v4825; shift_adder #(18, 13, 1, 1, 19, 4, 0) op_4825 (v3155[17:0], v2879[12:0], v4825[18:0]); // 4.0
    wire [20:0] v4826; shift_adder #(20, 13, 1, 1, 21, 7, 0) op_4826 (v3156[19:0], v3157[12:0], v4826[20:0]); // 4.0
    wire [19:0] v4827; shift_adder #(20, 15, 1, 1, 20, 3, 0) op_4827 (v3158[19:0], v3159[14:0], v4827[19:0]); // 4.0
    wire [23:0] v4828; shift_adder #(22, 23, 1, 1, 24, 0, 0) op_4828 (v3160[21:0], v3161[22:0], v4828[23:0]); // 4.0
    wire [20:0] v4829; shift_adder #(20, 20, 1, 1, 21, 0, 0) op_4829 (v3162[19:0], v3163[19:0], v4829[20:0]); // 4.0
    wire [18:0] v4830; shift_adder #(18, 16, 1, 1, 19, 2, 0) op_4830 (v3164[17:0], v3165[15:0], v4830[18:0]); // 4.0
    wire [22:0] v4831; shift_adder #(21, 20, 1, 1, 23, 2, 0) op_4831 (v3166[20:0], v3167[19:0], v4831[22:0]); // 4.0
    wire [23:0] v4832; shift_adder #(23, 16, 1, 1, 24, 8, 0) op_4832 (v3168[22:0], v3169[15:0], v4832[23:0]); // 4.0
    wire [24:0] v4833; shift_adder #(16, 24, 1, 1, 25, -7, 0) op_4833 (v3170[15:0], v3171[23:0], v4833[24:0]); // 4.0
    wire [28:0] v4834; shift_adder #(27, 20, 1, 1, 29, 8, 0) op_4834 (v3172[26:0], v3173[19:0], v4834[28:0]); // 4.0
    wire [25:0] v4835; shift_adder #(12, 26, 1, 1, 26, -12, 0) op_4835 (v3174[11:0], v3175[25:0], v4835[25:0]); // 4.0
    wire [23:0] v4836; shift_adder #(12, 23, 1, 1, 24, -12, 1) op_4836 (v1253[11:0], v3176[22:0], v4836[23:0]); // 4.0
    wire [15:0] v4837; shift_adder #(14, 13, 1, 1, 16, 2, 0) op_4837 (v2729[13:0], v3093[12:0], v4837[15:0]); // 4.0
    wire [20:0] v4838; shift_adder #(16, 20, 1, 1, 21, -4, 0) op_4838 (v3177[15:0], v3178[19:0], v4838[20:0]); // 4.0
    wire [17:0] v4839; shift_adder #(17, 17, 1, 1, 18, 0, 0) op_4839 (v3179[16:0], v3180[16:0], v4839[17:0]); // 4.0
    wire [19:0] v4840; shift_adder #(19, 17, 1, 1, 20, 2, 0) op_4840 (v2670[18:0], v3181[16:0], v4840[19:0]); // 4.0
    wire [23:0] v4841; shift_adder #(22, 23, 1, 1, 24, 1, 0) op_4841 (v3182[21:0], v3183[22:0], v4841[23:0]); // 4.0
    wire [26:0] v4842; shift_adder #(12, 27, 1, 1, 27, -9, 1) op_4842 (v151[11:0], v3184[26:0], v4842[26:0]); // 4.0
    wire [28:0] v4843; shift_adder #(23, 29, 1, 1, 29, -5, 0) op_4843 (v2666[22:0], v3185[28:0], v4843[28:0]); // 4.0
    wire [17:0] v4844; shift_adder #(15, 18, 1, 1, 18, 0, 0) op_4844 (v3186[14:0], v3187[17:0], v4844[17:0]); // 4.0
    wire [30:0] v4845; shift_adder #(11, 31, 1, 1, 31, -9, 1) op_4845 (v177[10:0], v3189[30:0], v4845[30:0]); // 4.0
    wire [27:0] v4846; shift_adder #(23, 28, 1, 1, 28, -4, 0) op_4846 (v3190[22:0], v3191[27:0], v4846[27:0]); // 4.0
    wire [38:0] v4847; shift_adder #(38, 34, 1, 1, 39, 4, 0) op_4847 (v3192[37:0], v3193[33:0], v4847[38:0]); // 4.0
    wire [35:0] v4848; shift_adder #(14, 13, 1, 1, 36, 23, 1) op_4848 (v3194[13:0], v1601[12:0], v4848[35:0]); // 4.0
    wire [24:0] v4849; shift_adder #(24, 16, 1, 1, 25, 9, 0) op_4849 (v3195[23:0], v3196[15:0], v4849[24:0]); // 4.0
    wire [39:0] v4850; shift_adder #(39, 22, 1, 1, 40, 18, 0) op_4850 (v3197[38:0], v3198[21:0], v4850[39:0]); // 4.0
    wire [17:0] v4851; shift_adder #(18, 14, 1, 1, 18, 2, 0) op_4851 (v3199[17:0], v3200[13:0], v4851[17:0]); // 4.0
    wire [16:0] v4852; shift_adder #(15, 15, 1, 1, 17, 1, 0) op_4852 (v3201[14:0], v3202[14:0], v4852[16:0]); // 4.0
    wire [17:0] v4853; shift_adder #(13, 18, 1, 1, 18, -2, 0) op_4853 (v3107[12:0], v3203[17:0], v4853[17:0]); // 4.0
    wire [15:0] v4854; shift_adder #(14, 16, 1, 1, 16, 0, 0) op_4854 (v3204[13:0], v3205[15:0], v4854[15:0]); // 4.0
    wire [19:0] v4855; shift_adder #(14, 20, 1, 1, 20, -3, 0) op_4855 (v3206[13:0], v2759[19:0], v4855[19:0]); // 4.0
    wire [15:0] v4856; shift_adder #(8, 16, 1, 1, 16, -3, 0) op_4856 (v69[7:0], v3207[15:0], v4856[15:0]); // 4.0
    wire [19:0] v4857; shift_adder #(18, 18, 1, 1, 20, -1, 0) op_4857 (v3208[17:0], v3209[17:0], v4857[19:0]); // 4.0
    wire [25:0] v4858; shift_adder #(23, 26, 1, 1, 26, -1, 0) op_4858 (v3210[22:0], v3211[25:0], v4858[25:0]); // 4.0
    wire [25:0] v4859; shift_adder #(24, 18, 1, 1, 26, 8, 0) op_4859 (v3212[23:0], v3213[17:0], v4859[25:0]); // 4.0
    wire [29:0] v4860; shift_adder #(25, 28, 1, 1, 30, -4, 0) op_4860 (v3214[24:0], v3215[27:0], v4860[29:0]); // 4.0
    wire [18:0] v4861; shift_adder #(12, 19, 1, 1, 19, 0, 1) op_4861 (v383[11:0], v3216[18:0], v4861[18:0]); // 4.0
    wire [23:0] v4862; shift_adder #(19, 24, 1, 1, 24, -3, 0) op_4862 (v3217[18:0], v3212[23:0], v4862[23:0]); // 4.0
    wire [20:0] v4863; shift_adder #(14, 20, 1, 1, 21, -5, 0) op_4863 (v3218[13:0], v3219[19:0], v4863[20:0]); // 4.0
    wire [19:0] v4864; shift_adder #(19, 19, 1, 1, 20, -1, 0) op_4864 (v3220[18:0], v3221[18:0], v4864[19:0]); // 4.0
    wire [21:0] v4865; shift_adder #(11, 22, 1, 1, 22, -6, 0) op_4865 (v168[10:0], v3222[21:0], v4865[21:0]); // 4.0
    wire [21:0] v4866; shift_adder #(21, 18, 1, 1, 22, 3, 0) op_4866 (v3223[20:0], v3068[17:0], v4866[21:0]); // 4.0
    wire [22:0] v4867; shift_adder #(22, 15, 1, 1, 23, 6, 0) op_4867 (v3224[21:0], v3225[14:0], v4867[22:0]); // 4.0
    wire [23:0] v4868; shift_adder #(16, 24, 1, 1, 24, -7, 0) op_4868 (v3165[15:0], v3195[23:0], v4868[23:0]); // 4.0
    wire [17:0] v4869; shift_adder #(11, 17, 1, 1, 18, -6, 1) op_4869 (v303[10:0], v3226[16:0], v4869[17:0]); // 4.0
    wire [31:0] v4870; shift_adder #(11, 24, 1, 1, 32, -21, 0) op_4870 (v284[10:0], v3227[23:0], v4870[31:0]); // 4.0
    wire [25:0] v4871; shift_adder #(18, 25, 1, 1, 26, -6, 0) op_4871 (v3228[17:0], v3229[24:0], v4871[25:0]); // 4.0
    wire [23:0] v4872; shift_adder #(22, 23, 1, 1, 24, -1, 0) op_4872 (v2682[21:0], v3230[22:0], v4872[23:0]); // 4.0
    wire [25:0] v4873; shift_adder #(25, 17, 1, 1, 26, 8, 0) op_4873 (v2715[24:0], v3231[16:0], v4873[25:0]); // 4.0
    wire [14:0] v4874; shift_adder #(14, 13, 1, 1, 15, 2, 0) op_4874 (v3232[13:0], v2522[12:0], v4874[14:0]); // 4.0
    wire [18:0] v4875; shift_adder #(16, 14, 1, 1, 19, 4, 0) op_4875 (v3233[15:0], v3234[13:0], v4875[18:0]); // 4.0
    wire [26:0] v4876; shift_adder #(26, 14, 1, 1, 27, 12, 0) op_4876 (v3235[25:0], v3236[13:0], v4876[26:0]); // 4.0
    wire [20:0] v4877; shift_adder #(20, 19, 1, 1, 21, 1, 0) op_4877 (v3237[19:0], v3238[18:0], v4877[20:0]); // 4.0
    wire [37:0] v4878; shift_adder #(14, 37, 1, 1, 38, -23, 0) op_4878 (v2692[13:0], v3239[36:0], v4878[37:0]); // 4.0
    wire [30:0] v4879; shift_adder #(29, 25, 1, 1, 31, 5, 0) op_4879 (v3240[28:0], v3241[24:0], v4879[30:0]); // 4.0
    wire [25:0] v4880; shift_adder #(25, 19, 1, 1, 26, 7, 0) op_4880 (v3242[24:0], v3243[18:0], v4880[25:0]); // 4.0
    wire [23:0] v4881; shift_adder #(22, 16, 1, 1, 24, 7, 0) op_4881 (v3244[21:0], v2787[15:0], v4881[23:0]); // 4.0
    wire [33:0] v4882; shift_adder #(22, 33, 1, 1, 34, -11, 0) op_4882 (v3245[21:0], v3246[32:0], v4882[33:0]); // 4.0
    wire [29:0] v4883; shift_adder #(23, 28, 1, 1, 30, -6, 0) op_4883 (v3247[22:0], v3248[27:0], v4883[29:0]); // 4.0
    wire [31:0] v4884; shift_adder #(31, 25, 1, 1, 32, 6, 0) op_4884 (v2539[30:0], v3249[24:0], v4884[31:0]); // 4.0
    wire [28:0] v4885; shift_adder #(13, 29, 1, 1, 29, -13, 1) op_4885 (v1660[12:0], v3250[28:0], v4885[28:0]); // 4.0
    wire [25:0] v4886; shift_adder #(26, 14, 1, 1, 26, 10, 0) op_4886 (v3251[25:0], v3252[13:0], v4886[25:0]); // 4.0
    wire [27:0] v4887; shift_adder #(28, 23, 1, 1, 28, 3, 0) op_4887 (v3253[27:0], v3254[22:0], v4887[27:0]); // 4.0
    wire [19:0] v4888; shift_adder #(17, 20, 1, 1, 20, -1, 0) op_4888 (v2559[16:0], v3255[19:0], v4888[19:0]); // 4.0
    wire [30:0] v4889; shift_adder #(22, 30, 1, 1, 31, -8, 0) op_4889 (v3245[21:0], v3256[29:0], v4889[30:0]); // 4.0
    wire [23:0] v4890; shift_adder #(23, 13, 1, 1, 24, 8, 0) op_4890 (v3257[22:0], v3258[12:0], v4890[23:0]); // 4.0
    wire [23:0] v4891; shift_adder #(16, 23, 1, 1, 24, -6, 0) op_4891 (v3259[15:0], v3260[22:0], v4891[23:0]); // 4.0
    wire [22:0] v4892; shift_adder #(22, 20, 1, 1, 23, 2, 0) op_4892 (v3261[21:0], v3262[19:0], v4892[22:0]); // 4.0
    wire [21:0] v4893; shift_adder #(22, 19, 1, 1, 22, 0, 0) op_4893 (v3263[21:0], v2516[18:0], v4893[21:0]); // 4.0
    wire [19:0] v4894; shift_adder #(19, 17, 1, 1, 20, 2, 0) op_4894 (v3264[18:0], v3265[16:0], v4894[19:0]); // 4.0
    wire [19:0] v4895; shift_adder #(14, 18, 1, 1, 20, -5, 0) op_4895 (v3266[13:0], v3267[17:0], v4895[19:0]); // 4.0
    wire [20:0] v4896; shift_adder #(16, 15, 1, 1, 21, 6, 0) op_4896 (v2513[15:0], v3268[14:0], v4896[20:0]); // 4.0
    wire [21:0] v4897; shift_adder #(16, 21, 1, 1, 22, -4, 0) op_4897 (v3269[15:0], v3270[20:0], v4897[21:0]); // 4.0
    wire [18:0] v4898; shift_adder #(19, 17, 1, 1, 19, 1, 0) op_4898 (v3271[18:0], v3272[16:0], v4898[18:0]); // 4.0
    wire [15:0] v4899; shift_adder #(14, 14, 1, 1, 16, 2, 0) op_4899 (v3273[13:0], v3002[13:0], v4899[15:0]); // 4.0
    wire [21:0] v4900; shift_adder #(17, 21, 1, 1, 22, -3, 0) op_4900 (v3274[16:0], v3275[20:0], v4900[21:0]); // 4.0
    wire [17:0] v4901; shift_adder #(10, 18, 1, 1, 18, -5, 1) op_4901 (v520[9:0], v3276[17:0], v4901[17:0]); // 4.0
    wire [24:0] v4902; shift_adder #(22, 23, 1, 1, 25, 1, 0) op_4902 (v3277[21:0], v3278[22:0], v4902[24:0]); // 4.0
    wire [19:0] v4903; shift_adder #(8, 17, 1, 1, 20, -11, 0) op_4903 (v68[7:0], v3279[16:0], v4903[19:0]); // 4.0
    wire [34:0] v4904; shift_adder #(19, 33, 1, 1, 35, -16, 0) op_4904 (v3280[18:0], v3281[32:0], v4904[34:0]); // 4.0
    wire [18:0] v4905; shift_adder #(18, 15, 1, 1, 19, 3, 0) op_4905 (v2727[17:0], v3016[14:0], v4905[18:0]); // 4.0
    wire [29:0] v4906; shift_adder #(29, 13, 1, 1, 30, 16, 0) op_4906 (v3282[28:0], v3283[12:0], v4906[29:0]); // 4.0
    wire [18:0] v4907; shift_adder #(18, 14, 1, 1, 19, 4, 0) op_4907 (v3284[17:0], v2776[13:0], v4907[18:0]); // 4.0
    wire [32:0] v4908; shift_adder #(18, 32, 1, 1, 33, -14, 0) op_4908 (v3285[17:0], v3286[31:0], v4908[32:0]); // 4.0
    wire [22:0] v4909; shift_adder #(20, 17, 1, 1, 23, 6, 0) op_4909 (v3287[19:0], v3288[16:0], v4909[22:0]); // 4.0
    wire [25:0] v4910; shift_adder #(20, 26, 1, 1, 26, -4, 0) op_4910 (v3289[19:0], v3043[25:0], v4910[25:0]); // 4.0
    wire [28:0] v4911; shift_adder #(20, 28, 1, 1, 29, -8, 0) op_4911 (v3290[19:0], v3291[27:0], v4911[28:0]); // 4.0
    wire [27:0] v4912; shift_adder #(20, 28, 1, 1, 28, -7, 0) op_4912 (v3292[19:0], v3293[27:0], v4912[27:0]); // 4.0
    wire [21:0] v4913; shift_adder #(20, 19, 1, 1, 22, 2, 0) op_4913 (v3287[19:0], v3294[18:0], v4913[21:0]); // 4.0
    wire [35:0] v4914; shift_adder #(33, 35, 1, 1, 36, -3, 0) op_4914 (v3295[32:0], v3296[34:0], v4914[35:0]); // 4.0
    wire [32:0] v4915; shift_adder #(32, 22, 1, 1, 33, 10, 0) op_4915 (v3076[31:0], v2770[21:0], v4915[32:0]); // 4.0
    wire [38:0] v4916; shift_adder #(17, 16, 1, 1, 39, 23, 1) op_4916 (v3297[16:0], v1275[15:0], v4916[38:0]); // 4.0
    wire [33:0] v4917; shift_adder #(34, 33, 1, 1, 34, 0, 0) op_4917 (v3298[33:0], v3299[32:0], v4917[33:0]); // 4.0
    wire [35:0] v4918; shift_adder #(29, 15, 1, 1, 36, -7, 1) op_4918 (v3300[28:0], v3301[14:0], v4918[35:0]); // 4.0
    wire [36:0] v4919; shift_adder #(12, 36, 1, 1, 37, -24, 0) op_4919 (v3302[11:0], v3303[35:0], v4919[36:0]); // 4.0
    wire [22:0] v4920; shift_adder #(23, 16, 1, 1, 23, 4, 0) op_4920 (v3304[22:0], v3305[15:0], v4920[22:0]); // 4.0
    wire [19:0] v4921; shift_adder #(18, 19, 1, 1, 20, -1, 0) op_4921 (v3018[17:0], v3306[18:0], v4921[19:0]); // 4.0
    wire [17:0] v4922; shift_adder #(11, 16, 1, 1, 18, -7, 0) op_4922 (v341[10:0], v3307[15:0], v4922[17:0]); // 4.0
    wire [17:0] v4923; shift_adder #(15, 16, 1, 1, 18, 1, 0) op_4923 (v3308[14:0], v3309[15:0], v4923[17:0]); // 4.0
    wire [21:0] v4924; shift_adder #(17, 22, 1, 1, 22, -4, 0) op_4924 (v2696[16:0], v3310[21:0], v4924[21:0]); // 4.0
    wire [32:0] v4925; shift_adder #(32, 16, 1, 1, 33, 16, 0) op_4925 (v3311[31:0], v3312[15:0], v4925[32:0]); // 4.0
    wire [28:0] v4926; shift_adder #(22, 28, 1, 1, 29, -6, 0) op_4926 (v3313[21:0], v3314[27:0], v4926[28:0]); // 4.0
    wire [30:0] v4927; shift_adder #(31, 29, 1, 1, 31, 1, 0) op_4927 (v2782[30:0], v3315[28:0], v4927[30:0]); // 4.0
    wire [30:0] v4928; shift_adder #(31, 15, 1, 1, 31, 15, 0) op_4928 (v3316[30:0], v2721[14:0], v4928[30:0]); // 4.0
    wire [28:0] v4929; shift_adder #(27, 20, 1, 1, 29, 8, 0) op_4929 (v3317[26:0], v3318[19:0], v4929[28:0]); // 4.0
    wire [23:0] v4930; shift_adder #(19, 23, 1, 1, 24, -4, 0) op_4930 (v3319[18:0], v3320[22:0], v4930[23:0]); // 4.0
    wire [24:0] v4931; shift_adder #(22, 25, 1, 1, 25, -2, 0) op_4931 (v3321[21:0], v3322[24:0], v4931[24:0]); // 4.0
    wire [26:0] v4932; shift_adder #(20, 26, 1, 1, 27, -5, 0) op_4932 (v3323[19:0], v3324[25:0], v4932[26:0]); // 4.0
    wire [28:0] v4933; shift_adder #(28, 14, 1, 1, 29, 13, 0) op_4933 (v3325[27:0], v3326[13:0], v4933[28:0]); // 4.0
    wire [27:0] v4934; shift_adder #(23, 28, 1, 1, 28, -4, 0) op_4934 (v3327[22:0], v3328[27:0], v4934[27:0]); // 4.0
    wire [22:0] v4935; shift_adder #(18, 22, 1, 1, 23, -3, 0) op_4935 (v3329[17:0], v3330[21:0], v4935[22:0]); // 4.0
    wire [21:0] v4936; shift_adder #(20, 21, 1, 1, 22, -1, 0) op_4936 (v3059[19:0], v3331[20:0], v4936[21:0]); // 4.0
    wire [19:0] v4937; shift_adder #(20, 16, 1, 1, 20, 2, 0) op_4937 (v3332[19:0], v3333[15:0], v4937[19:0]); // 4.0
    wire [24:0] v4938; shift_adder #(25, 18, 1, 1, 25, 3, 1) op_4938 (v791[24:0], v2761[17:0], v4938[24:0]); // 4.0
    wire [19:0] v4939; shift_adder #(15, 20, 1, 1, 20, -3, 0) op_4939 (v3334[14:0], v3335[19:0], v4939[19:0]); // 4.0
    wire [24:0] v4940; shift_adder #(23, 16, 1, 1, 25, 8, 0) op_4940 (v3336[22:0], v3337[15:0], v4940[24:0]); // 4.0
    wire [22:0] v4941; shift_adder #(20, 23, 1, 1, 23, -1, 0) op_4941 (v3338[19:0], v3339[22:0], v4941[22:0]); // 4.0
    wire [31:0] v4942; shift_adder #(31, 28, 1, 1, 32, 3, 0) op_4942 (v3340[30:0], v2926[27:0], v4942[31:0]); // 4.0
    wire [32:0] v4943; shift_adder #(33, 24, 1, 1, 33, 8, 0) op_4943 (v3295[32:0], v3341[23:0], v4943[32:0]); // 4.0
    wire [31:0] v4944; shift_adder #(24, 30, 1, 1, 32, -7, 0) op_4944 (v3342[23:0], v3343[29:0], v4944[31:0]); // 4.0
    wire [22:0] v4945; shift_adder #(22, 15, 1, 1, 23, 7, 0) op_4945 (v3344[21:0], v3345[14:0], v4945[22:0]); // 4.0
    wire [28:0] v4946; shift_adder #(13, 29, 1, 1, 29, -13, 0) op_4946 (v3119[12:0], v2798[28:0], v4946[28:0]); // 4.0
    wire [25:0] v4947; shift_adder #(11, 15, 1, 1, 26, 11, 1) op_4947 (v134[10:0], v3346[14:0], v4947[25:0]); // 4.0
    wire [30:0] v4948; shift_adder #(22, 30, 1, 1, 31, -8, 0) op_4948 (v3347[21:0], v3348[29:0], v4948[30:0]); // 4.0
    wire [27:0] v4949; shift_adder #(26, 25, 1, 1, 28, 2, 0) op_4949 (v3349[25:0], v3350[24:0], v4949[27:0]); // 4.0
    wire [22:0] v4950; shift_adder #(21, 21, 1, 1, 23, 1, 0) op_4950 (v2885[20:0], v2909[20:0], v4950[22:0]); // 4.0
    wire [22:0] v4951; shift_adder #(18, 22, 1, 1, 23, -4, 0) op_4951 (v3164[17:0], v3351[21:0], v4951[22:0]); // 4.0
    wire [19:0] v4952; shift_adder #(20, 17, 1, 1, 20, 2, 0) op_4952 (v3352[19:0], v3353[16:0], v4952[19:0]); // 4.0
    wire [25:0] v4953; shift_adder #(15, 24, 1, 1, 26, -10, 0) op_4953 (v3354[14:0], v3355[23:0], v4953[25:0]); // 4.0
    wire [15:0] v4954; shift_adder #(13, 15, 1, 1, 16, -1, 0) op_4954 (v3356[12:0], v3357[14:0], v4954[15:0]); // 4.0
    wire [22:0] v4955; shift_adder #(23, 15, 1, 1, 23, 7, 0) op_4955 (v3183[22:0], v3358[14:0], v4955[22:0]); // 4.0
    wire [24:0] v4956; shift_adder #(24, 15, 1, 1, 25, 10, 0) op_4956 (v3359[23:0], v2987[14:0], v4956[24:0]); // 4.0
    wire [23:0] v4957; shift_adder #(23, 18, 1, 1, 24, 5, 0) op_4957 (v3360[22:0], v3361[17:0], v4957[23:0]); // 4.0
    wire [32:0] v4958; shift_adder #(8, 33, 1, 1, 33, -10, 1) op_4958 (v77[7:0], v3362[32:0], v4958[32:0]); // 4.0
    wire [28:0] v4959; shift_adder #(14, 13, 1, 1, 29, 16, 0) op_4959 (v1378[13:0], v3363[12:0], v4959[28:0]); // 4.0
    wire [29:0] v4960; shift_adder #(24, 30, 1, 1, 30, -5, 0) op_4960 (v3364[23:0], v3365[29:0], v4960[29:0]); // 4.0
    wire [17:0] v4961; shift_adder #(15, 16, 1, 1, 18, 2, 0) op_4961 (v3366[14:0], v3367[15:0], v4961[17:0]); // 4.0
    wire [18:0] v4962; shift_adder #(17, 14, 1, 1, 19, 4, 0) op_4962 (v3368[16:0], v3369[13:0], v4962[18:0]); // 4.0
    wire [35:0] v4963; shift_adder #(35, 19, 1, 1, 36, 16, 0) op_4963 (v3370[34:0], v3371[18:0], v4963[35:0]); // 4.0
    wire [29:0] v4964; shift_adder #(28, 16, 1, 1, 30, 13, 0) op_4964 (v3372[27:0], v3373[15:0], v4964[29:0]); // 4.0
    wire [33:0] v4965; shift_adder #(33, 16, 1, 1, 34, 18, 0) op_4965 (v3374[32:0], v3375[15:0], v4965[33:0]); // 4.0
    wire [33:0] v4966; shift_adder #(19, 34, 1, 1, 34, -13, 0) op_4966 (v3376[18:0], v3377[33:0], v4966[33:0]); // 4.0
    wire [37:0] v4967; shift_adder #(14, 28, 1, 1, 38, 10, 1) op_4967 (v3378[13:0], v1777[27:0], v4967[37:0]); // 4.0
    wire [24:0] v4968; shift_adder #(13, 24, 1, 1, 25, -11, 0) op_4968 (v2929[12:0], v3379[23:0], v4968[24:0]); // 4.0
    wire [34:0] v4969; shift_adder #(25, 34, 1, 1, 35, -9, 0) op_4969 (v3380[24:0], v3381[33:0], v4969[34:0]); // 4.0
    wire [18:0] v4970; shift_adder #(14, 18, 1, 1, 19, -4, 0) op_4970 (v3382[13:0], v3383[17:0], v4970[18:0]); // 4.0
    wire [37:0] v4971; shift_adder #(15, 37, 1, 1, 38, -23, 0) op_4971 (v3384[14:0], v3385[36:0], v4971[37:0]); // 4.0
    wire [16:0] v4972; shift_adder #(15, 15, 1, 1, 17, -2, 0) op_4972 (v3386[14:0], v3387[14:0], v4972[16:0]); // 4.0
    wire [19:0] v4973; shift_adder #(14, 20, 1, 1, 20, -5, 0) op_4973 (v2788[13:0], v3388[19:0], v4973[19:0]); // 4.0
    wire [21:0] v4974; shift_adder #(15, 21, 1, 1, 22, -6, 0) op_4974 (v3389[14:0], v3390[20:0], v4974[21:0]); // 4.0
    wire [21:0] v4975; shift_adder #(21, 20, 1, 1, 22, 0, 0) op_4975 (v3391[20:0], v3392[19:0], v4975[21:0]); // 4.0
    wire [25:0] v4976; shift_adder #(26, 21, 1, 1, 26, 3, 0) op_4976 (v3393[25:0], v3394[20:0], v4976[25:0]); // 4.0
    wire [16:0] v4977; shift_adder #(14, 16, 1, 1, 17, -3, 0) op_4977 (v3395[13:0], v3396[15:0], v4977[16:0]); // 4.0
    wire [17:0] v4978; shift_adder #(17, 17, 1, 1, 18, 0, 0) op_4978 (v3397[16:0], v3398[16:0], v4978[17:0]); // 4.0
    wire [18:0] v4979; shift_adder #(17, 16, 1, 1, 19, 2, 0) op_4979 (v3353[16:0], v3399[15:0], v4979[18:0]); // 4.0
    wire [24:0] v4980; shift_adder #(23, 24, 1, 1, 25, -1, 0) op_4980 (v3400[22:0], v3401[23:0], v4980[24:0]); // 4.0
    wire [21:0] v4981; shift_adder #(19, 21, 1, 1, 22, -1, 0) op_4981 (v3402[18:0], v3403[20:0], v4981[21:0]); // 4.0
    wire [19:0] v4982; shift_adder #(13, 19, 1, 1, 20, -6, 0) op_4982 (v2612[12:0], v3404[18:0], v4982[19:0]); // 4.0
    wire [17:0] v4983; shift_adder #(16, 18, 1, 1, 18, -1, 0) op_4983 (v3405[15:0], v3406[17:0], v4983[17:0]); // 4.0
    wire [29:0] v4984; shift_adder #(17, 30, 1, 1, 30, -12, 0) op_4984 (v3407[16:0], v3408[29:0], v4984[29:0]); // 4.0
    wire [27:0] v4985; shift_adder #(20, 27, 1, 1, 28, -6, 0) op_4985 (v3066[19:0], v3409[26:0], v4985[27:0]); // 4.0
    wire [26:0] v4986; shift_adder #(15, 20, 1, 1, 27, 7, 0) op_4986 (v253[14:0], v3410[19:0], v4986[26:0]); // 4.0
    wire [18:0] v4987; shift_adder #(16, 18, 1, 1, 19, -1, 0) op_4987 (v2863[15:0], v3411[17:0], v4987[18:0]); // 4.0
    wire [22:0] v4988; shift_adder #(21, 19, 1, 1, 23, 3, 0) op_4988 (v3412[20:0], v3413[18:0], v4988[22:0]); // 4.0
    wire [27:0] v4989; shift_adder #(11, 25, 1, 1, 28, 3, 1) op_4989 (v846[10:0], v3414[24:0], v4989[27:0]); // 4.0
    wire [28:0] v4990; shift_adder #(28, 19, 1, 1, 29, 10, 0) op_4990 (v3415[27:0], v3416[18:0], v4990[28:0]); // 4.0
    wire [35:0] v4991; shift_adder #(12, 36, 1, 1, 36, -23, 0) op_4991 (v3417[11:0], v3418[35:0], v4991[35:0]); // 4.0
    wire [18:0] v4992; shift_adder #(15, 19, 1, 1, 19, -2, 0) op_4992 (v3419[14:0], v2773[18:0], v4992[18:0]); // 4.0
    wire [16:0] v4993; shift_adder #(16, 13, 1, 1, 17, 3, 0) op_4993 (v3420[15:0], v3421[12:0], v4993[16:0]); // 4.0
    wire [33:0] v4994; shift_adder #(19, 33, 1, 1, 34, -14, 0) op_4994 (v3422[18:0], v3423[32:0], v4994[33:0]); // 4.0
    wire [22:0] v4995; shift_adder #(22, 19, 1, 1, 23, 3, 0) op_4995 (v3424[21:0], v3425[18:0], v4995[22:0]); // 4.0
    wire [29:0] v4996; shift_adder #(20, 29, 1, 1, 30, -9, 0) op_4996 (v2590[19:0], v3426[28:0], v4996[29:0]); // 4.0
    wire [38:0] v4997; shift_adder #(18, 14, 1, 1, 39, -21, 1) op_4997 (v3427[17:0], v3428[13:0], v4997[38:0]); // 4.0
    wire [25:0] v4998; shift_adder #(25, 23, 1, 1, 26, 1, 0) op_4998 (v3133[24:0], v3429[22:0], v4998[25:0]); // 4.0
    wire [16:0] v4999; shift_adder #(15, 15, 1, 1, 17, 1, 0) op_4999 (v3430[14:0], v2555[14:0], v4999[16:0]); // 4.0
    wire [22:0] v5000; shift_adder #(23, 17, 1, 1, 23, 4, 0) op_5000 (v3431[22:0], v3432[16:0], v5000[22:0]); // 4.0
    wire [18:0] v5001; shift_adder #(17, 15, 1, 1, 19, 3, 0) op_5001 (v2529[16:0], v3433[14:0], v5001[18:0]); // 4.0
    wire [19:0] v5002; shift_adder #(20, 18, 1, 1, 20, 0, 0) op_5002 (v3434[19:0], v3435[17:0], v5002[19:0]); // 4.0
    wire [17:0] v5003; shift_adder #(16, 17, 1, 1, 18, -1, 0) op_5003 (v3436[15:0], v3279[16:0], v5003[17:0]); // 4.0
    wire [18:0] v5004; shift_adder #(16, 16, 1, 1, 19, -2, 0) op_5004 (v3437[15:0], v3438[15:0], v5004[18:0]); // 4.0
    wire [16:0] v5005; shift_adder #(16, 15, 1, 1, 17, 0, 0) op_5005 (v3439[15:0], v3440[14:0], v5005[16:0]); // 4.0
    wire [24:0] v5006; shift_adder #(24, 15, 1, 1, 25, 8, 0) op_5006 (v3441[23:0], v3442[14:0], v5006[24:0]); // 4.0
    wire [25:0] v5007; shift_adder #(15, 26, 1, 1, 26, -10, 0) op_5007 (v3443[14:0], v3444[25:0], v5007[25:0]); // 4.0
    wire [17:0] v5008; shift_adder #(16, 16, 1, 1, 18, -1, 0) op_5008 (v3445[15:0], v3446[15:0], v5008[17:0]); // 4.0
    wire [25:0] v5009; shift_adder #(26, 20, 1, 1, 26, 4, 0) op_5009 (v3447[25:0], v3448[19:0], v5009[25:0]); // 4.0
    wire [23:0] v5010; shift_adder #(14, 22, 1, 1, 24, -10, 0) op_5010 (v2908[13:0], v3449[21:0], v5010[23:0]); // 4.0
    wire [23:0] v5011; shift_adder #(11, 24, 1, 1, 24, -3, 0) op_5011 (v133[10:0], v3450[23:0], v5011[23:0]); // 4.0
    wire [27:0] v5012; shift_adder #(27, 24, 1, 1, 28, 3, 0) op_5012 (v3077[26:0], v3451[23:0], v5012[27:0]); // 4.0
    wire [18:0] v5013; shift_adder #(16, 18, 1, 1, 19, -2, 0) op_5013 (v3452[15:0], v3285[17:0], v5013[18:0]); // 4.0
    wire [29:0] v5014; shift_adder #(30, 26, 1, 1, 30, 1, 0) op_5014 (v2681[29:0], v3453[25:0], v5014[29:0]); // 4.0
    wire [24:0] v5015; shift_adder #(25, 18, 1, 1, 25, 5, 0) op_5015 (v3454[24:0], v3455[17:0], v5015[24:0]); // 4.0
    wire [25:0] v5016; shift_adder #(25, 25, 1, 1, 26, -1, 0) op_5016 (v3456[24:0], v3457[24:0], v5016[25:0]); // 4.0
    wire [19:0] v5017; shift_adder #(19, 14, 1, 1, 20, 5, 0) op_5017 (v3458[18:0], v3459[13:0], v5017[19:0]); // 4.0
    wire [25:0] v5018; shift_adder #(21, 26, 1, 1, 26, -3, 0) op_5018 (v3460[20:0], v3461[25:0], v5018[25:0]); // 4.0
    wire [19:0] v5019; shift_adder #(18, 19, 1, 1, 20, 1, 0) op_5019 (v3462[17:0], v3463[18:0], v5019[19:0]); // 4.0
    wire [17:0] v5020; shift_adder #(8, 18, 1, 1, 18, -1, 1) op_5020 (v66[7:0], v3464[17:0], v5020[17:0]); // 4.0
    wire [21:0] v5021; shift_adder #(20, 19, 1, 1, 22, 2, 0) op_5021 (v3465[19:0], v3466[18:0], v5021[21:0]); // 4.0
    wire [25:0] v5022; shift_adder #(17, 26, 1, 1, 26, -7, 0) op_5022 (v3467[16:0], v3468[25:0], v5022[25:0]); // 4.0
    wire [20:0] v5023; shift_adder #(20, 13, 1, 1, 21, 8, 0) op_5023 (v3469[19:0], v3363[12:0], v5023[20:0]); // 4.0
    wire [19:0] v5024; shift_adder #(19, 15, 1, 1, 20, 4, 0) op_5024 (v3470[18:0], v2709[14:0], v5024[19:0]); // 4.0
    wire [19:0] v5025; shift_adder #(19, 20, 1, 1, 20, 0, 0) op_5025 (v2658[18:0], v3448[19:0], v5025[19:0]); // 4.0
    wire [18:0] v5026; shift_adder #(17, 18, 1, 1, 19, -1, 0) op_5026 (v3471[16:0], v3131[17:0], v5026[18:0]); // 4.0
    wire [23:0] v5027; shift_adder #(15, 24, 1, 1, 24, -7, 0) op_5027 (v2914[14:0], v2514[23:0], v5027[23:0]); // 4.0
    wire [28:0] v5028; shift_adder #(28, 26, 1, 1, 29, 2, 0) op_5028 (v3472[27:0], v3473[25:0], v5028[28:0]); // 4.0
    wire [27:0] v5029; shift_adder #(27, 20, 1, 1, 28, 6, 0) op_5029 (v3474[26:0], v3392[19:0], v5029[27:0]); // 4.0
    wire [26:0] v5030; shift_adder #(26, 22, 1, 1, 27, 4, 0) op_5030 (v3251[25:0], v3475[21:0], v5030[26:0]); // 4.0
    wire [26:0] v5031; shift_adder #(24, 23, 1, 1, 27, 4, 0) op_5031 (v3476[23:0], v2616[22:0], v5031[26:0]); // 4.0
    wire [19:0] v5032; shift_adder #(19, 17, 1, 1, 20, 2, 0) op_5032 (v3477[18:0], v3353[16:0], v5032[19:0]); // 4.0
    wire [40:0] v5033; shift_adder #(20, 15, 1, 1, 41, 26, 1) op_5033 (v3478[19:0], v1861[14:0], v5033[40:0]); // 4.0
    wire [31:0] v5034; shift_adder #(8, 22, 1, 1, 32, -23, 0) op_5034 (v71[7:0], v3479[21:0], v5034[31:0]); // 4.0
    wire [14:0] v5035; shift_adder #(14, 13, 1, 1, 15, 1, 0) op_5035 (v3480[13:0], v3283[12:0], v5035[14:0]); // 4.0
    wire [27:0] v5036; shift_adder #(28, 14, 1, 1, 28, 12, 0) op_5036 (v3481[27:0], v3482[13:0], v5036[27:0]); // 4.0
    wire [18:0] v5037; shift_adder #(18, 18, 1, 1, 19, 0, 0) op_5037 (v3483[17:0], v2589[17:0], v5037[18:0]); // 4.0
    wire [16:0] v5038; shift_adder #(16, 16, 1, 1, 17, -1, 0) op_5038 (v3484[15:0], v3485[15:0], v5038[16:0]); // 4.0
    wire [18:0] v5039; shift_adder #(14, 18, 1, 1, 19, -4, 0) op_5039 (v2953[13:0], v3486[17:0], v5039[18:0]); // 4.0
    wire [19:0] v5040; shift_adder #(16, 15, 1, 1, 20, 4, 0) op_5040 (v3396[15:0], v2839[14:0], v5040[19:0]); // 4.0
    wire [20:0] v5041; shift_adder #(20, 17, 1, 1, 21, 3, 0) op_5041 (v3487[19:0], v3488[16:0], v5041[20:0]); // 4.0
    wire [19:0] v5042; shift_adder #(18, 19, 1, 1, 20, -1, 0) op_5042 (v3489[17:0], v3490[18:0], v5042[19:0]); // 4.0
    wire [34:0] v5043; shift_adder #(34, 34, 1, 1, 35, 0, 0) op_5043 (v3491[33:0], v3492[33:0], v5043[34:0]); // 4.0
    wire [37:0] v5044; shift_adder #(33, 37, 1, 1, 38, -3, 0) op_5044 (v3493[32:0], v3494[36:0], v5044[37:0]); // 4.0
    wire [16:0] v5045; shift_adder #(16, 14, 1, 1, 17, 2, 0) op_5045 (v3495[15:0], v3496[13:0], v5045[16:0]); // 4.0
    wire [16:0] v5046; shift_adder #(13, 16, 1, 1, 17, -3, 0) op_5046 (v2956[12:0], v3233[15:0], v5046[16:0]); // 4.0
    wire [33:0] v5047; shift_adder #(16, 33, 1, 1, 34, -17, 0) op_5047 (v3497[15:0], v3498[32:0], v5047[33:0]); // 4.0
    wire [14:0] v5048; shift_adder #(13, 14, 1, 1, 15, -2, 0) op_5048 (v3499[12:0], v3500[13:0], v5048[14:0]); // 4.0
    wire [22:0] v5049; shift_adder #(22, 22, 1, 1, 23, -1, 0) op_5049 (v3501[21:0], v3502[21:0], v5049[22:0]); // 4.0
    wire [23:0] v5050; shift_adder #(24, 20, 1, 1, 24, 2, 0) op_5050 (v3048[23:0], v3448[19:0], v5050[23:0]); // 4.0
    wire [31:0] v5051; shift_adder #(27, 30, 1, 1, 32, -4, 0) op_5051 (v3503[26:0], v3504[29:0], v5051[31:0]); // 4.0
    wire [28:0] v5052; shift_adder #(28, 13, 1, 1, 29, 15, 0) op_5052 (v3191[27:0], v3505[12:0], v5052[28:0]); // 4.0
    wire [26:0] v5053; shift_adder #(22, 26, 1, 1, 27, -5, 0) op_5053 (v2900[21:0], v3506[25:0], v5053[26:0]); // 4.0
    wire [22:0] v5054; shift_adder #(16, 22, 1, 1, 23, -6, 0) op_5054 (v3507[15:0], v3508[21:0], v5054[22:0]); // 4.0
    wire [28:0] v5055; shift_adder #(27, 24, 1, 1, 29, 4, 0) op_5055 (v3509[26:0], v3510[23:0], v5055[28:0]); // 4.0
    wire [30:0] v5056; shift_adder #(26, 29, 1, 1, 31, -4, 0) op_5056 (v3511[25:0], v3512[28:0], v5056[30:0]); // 4.0
    wire [19:0] v5057; shift_adder #(20, 14, 1, 1, 20, 4, 0) op_5057 (v3513[19:0], v3326[13:0], v5057[19:0]); // 4.0
    wire [18:0] v5058; shift_adder #(18, 14, 1, 1, 19, 4, 0) op_5058 (v3514[17:0], v3515[13:0], v5058[18:0]); // 4.0
    wire [24:0] v5059; shift_adder #(22, 25, 1, 1, 25, -1, 0) op_5059 (v3516[21:0], v3517[24:0], v5059[24:0]); // 4.0
    wire [22:0] v5060; shift_adder #(23, 17, 1, 1, 23, 4, 0) op_5060 (v3518[22:0], v3519[16:0], v5060[22:0]); // 4.0
    wire [23:0] v5061; shift_adder #(22, 19, 1, 1, 24, 4, 0) op_5061 (v3508[21:0], v3520[18:0], v5061[23:0]); // 4.0
    wire [16:0] v5062; shift_adder #(13, 16, 1, 1, 17, -3, 0) op_5062 (v2876[12:0], v3521[15:0], v5062[16:0]); // 4.0
    wire [21:0] v5063; shift_adder #(21, 19, 1, 1, 22, 2, 0) op_5063 (v3522[20:0], v2802[18:0], v5063[21:0]); // 4.0
    wire [18:0] v5064; shift_adder #(17, 18, 1, 1, 19, -1, 0) op_5064 (v2986[16:0], v3523[17:0], v5064[18:0]); // 4.0
    wire [20:0] v5065; shift_adder #(19, 13, 1, 1, 21, 7, 0) op_5065 (v2678[18:0], v3524[12:0], v5065[20:0]); // 4.0
    wire [22:0] v5066; shift_adder #(22, 22, 1, 1, 23, 1, 0) op_5066 (v3525[21:0], v3313[21:0], v5066[22:0]); // 4.0
    wire [23:0] v5067; shift_adder #(23, 22, 1, 1, 24, 2, 0) op_5067 (v3431[22:0], v3526[21:0], v5067[23:0]); // 4.0
    wire [32:0] v5068; shift_adder #(14, 33, 1, 1, 33, -15, 0) op_5068 (v3527[13:0], v3528[32:0], v5068[32:0]); // 4.0
    wire [23:0] v5069; shift_adder #(17, 23, 1, 1, 24, -5, 0) op_5069 (v3529[16:0], v3230[22:0], v5069[23:0]); // 4.0
    wire [22:0] v5070; shift_adder #(22, 20, 1, 1, 23, 3, 0) op_5070 (v3530[21:0], v3531[19:0], v5070[22:0]); // 4.0
    wire [32:0] v5071; shift_adder #(20, 33, 1, 1, 33, -10, 0) op_5071 (v3532[19:0], v3533[32:0], v5071[32:0]); // 4.0
    wire [24:0] v5072; shift_adder #(24, 23, 1, 1, 25, 1, 0) op_5072 (v3115[23:0], v3534[22:0], v5072[24:0]); // 4.0
    wire [24:0] v5073; shift_adder #(19, 24, 1, 1, 25, -5, 0) op_5073 (v3535[18:0], v3536[23:0], v5073[24:0]); // 4.0
    wire [38:0] v5074; shift_adder #(38, 20, 1, 1, 39, 19, 0) op_5074 (v3537[37:0], v3538[19:0], v5074[38:0]); // 4.0
    wire [40:0] v5075; shift_adder #(40, 16, 1, 1, 41, 25, 0) op_5075 (v3539[39:0], v3540[15:0], v5075[40:0]); // 4.0
    wire [18:0] v5076; shift_adder #(19, 13, 1, 1, 19, 4, 0) op_5076 (v3541[18:0], v3542[12:0], v5076[18:0]); // 4.0
    wire [25:0] v5077; shift_adder #(18, 25, 1, 1, 26, -7, 0) op_5077 (v3543[17:0], v2945[24:0], v5077[25:0]); // 4.0
    wire [16:0] v5078; shift_adder #(17, 14, 1, 1, 17, 2, 0) op_5078 (v3544[16:0], v3273[13:0], v5078[16:0]); // 4.0
    wire [17:0] v5079; shift_adder #(17, 16, 1, 1, 18, 0, 0) op_5079 (v3545[16:0], v3546[15:0], v5079[17:0]); // 4.0
    wire [19:0] v5080; shift_adder #(16, 20, 1, 1, 20, -3, 0) op_5080 (v3019[15:0], v3352[19:0], v5080[19:0]); // 4.0
    wire [15:0] v5081; shift_adder #(14, 14, 1, 1, 16, 2, 0) op_5081 (v3547[13:0], v3548[13:0], v5081[15:0]); // 4.0
    wire [17:0] v5082; shift_adder #(16, 14, 1, 1, 18, 4, 0) op_5082 (v3549[15:0], v3135[13:0], v5082[17:0]); // 4.0
    wire [35:0] v5083; shift_adder #(18, 36, 1, 1, 36, -17, 0) op_5083 (v3550[17:0], v3551[35:0], v5083[35:0]); // 4.0
    wire [35:0] v5084; shift_adder #(35, 21, 1, 1, 36, 14, 0) op_5084 (v2814[34:0], v3552[20:0], v5084[35:0]); // 4.0
    wire [21:0] v5085; shift_adder #(21, 20, 1, 1, 22, 1, 0) op_5085 (v3553[20:0], v3554[19:0], v5085[21:0]); // 4.0
    wire [18:0] v5086; shift_adder #(17, 16, 1, 1, 19, 2, 0) op_5086 (v2891[16:0], v3555[15:0], v5086[18:0]); // 4.0
    wire [15:0] v5087; shift_adder #(15, 14, 1, 1, 16, 0, 0) op_5087 (v3556[14:0], v3557[13:0], v5087[15:0]); // 4.0
    wire [31:0] v5088; shift_adder #(10, 31, 1, 1, 32, -21, 0) op_5088 (v130[9:0], v3558[30:0], v5088[31:0]); // 4.0
    wire [33:0] v5089; shift_adder #(28, 32, 1, 1, 34, -6, 0) op_5089 (v3559[27:0], v2812[31:0], v5089[33:0]); // 4.0
    wire [33:0] v5090; shift_adder #(24, 32, 1, 1, 34, -9, 0) op_5090 (v2881[23:0], v3560[31:0], v5090[33:0]); // 4.0
    wire [27:0] v5091; shift_adder #(27, 22, 1, 1, 28, 5, 0) op_5091 (v2724[26:0], v3561[21:0], v5091[27:0]); // 4.0
    wire [28:0] v5092; shift_adder #(18, 28, 1, 1, 29, -11, 0) op_5092 (v3562[17:0], v3563[27:0], v5092[28:0]); // 4.0
    wire [29:0] v5093; shift_adder #(28, 28, 1, 1, 30, 2, 0) op_5093 (v3564[27:0], v3565[27:0], v5093[29:0]); // 4.0
    wire [32:0] v5094; shift_adder #(21, 32, 1, 1, 33, -11, 0) op_5094 (v3566[20:0], v3567[31:0], v5094[32:0]); // 4.0
    wire [24:0] v5095; shift_adder #(24, 17, 1, 1, 25, 6, 0) op_5095 (v3568[23:0], v3569[16:0], v5095[24:0]); // 4.0
    wire [25:0] v5096; shift_adder #(25, 15, 1, 1, 26, 9, 0) op_5096 (v3570[24:0], v3571[14:0], v5096[25:0]); // 4.0
    wire [25:0] v5097; shift_adder #(26, 12, 1, 1, 26, 12, 0) op_5097 (v3099[25:0], v1068[11:0], v5097[25:0]); // 4.0
    wire [22:0] v5098; shift_adder #(16, 21, 1, 1, 23, -7, 0) op_5098 (v3572[15:0], v2628[20:0], v5098[22:0]); // 4.0
    wire [20:0] v5099; shift_adder #(20, 18, 1, 1, 21, 2, 0) op_5099 (v3573[19:0], v3574[17:0], v5099[20:0]); // 4.0
    wire [28:0] v5100; shift_adder #(11, 27, 1, 1, 29, 2, 1) op_5100 (v190[10:0], v3575[26:0], v5100[28:0]); // 4.0
    wire [21:0] v5101; shift_adder #(20, 20, 1, 1, 22, -2, 0) op_5101 (v3576[19:0], v3289[19:0], v5101[21:0]); // 4.0
    wire [25:0] v5102; shift_adder #(16, 26, 1, 1, 26, -6, 0) op_5102 (v3577[15:0], v3578[25:0], v5102[25:0]); // 4.0
    wire [29:0] v5103; shift_adder #(29, 24, 1, 1, 30, 5, 0) op_5103 (v3579[28:0], v3580[23:0], v5103[29:0]); // 4.0
    wire [29:0] v5104; shift_adder #(29, 15, 1, 1, 30, 13, 0) op_5104 (v3581[28:0], v3582[14:0], v5104[29:0]); // 4.0
    wire [25:0] v5105; shift_adder #(25, 14, 1, 1, 26, 10, 0) op_5105 (v3583[24:0], v3584[13:0], v5105[25:0]); // 4.0
    wire [19:0] v5106; shift_adder #(17, 19, 1, 1, 20, -2, 0) op_5106 (v3585[16:0], v3586[18:0], v5106[19:0]); // 4.0
    wire [25:0] v5107; shift_adder #(24, 15, 1, 1, 26, 10, 0) op_5107 (v2813[23:0], v3587[14:0], v5107[25:0]); // 4.0
    wire [15:0] v5108; shift_adder #(15, 13, 1, 1, 16, 1, 0) op_5108 (v3588[14:0], v2939[12:0], v5108[15:0]); // 4.0
    wire [20:0] v5109; shift_adder #(16, 21, 1, 1, 21, -2, 0) op_5109 (v3373[15:0], v3589[20:0], v5109[20:0]); // 4.0
    wire [22:0] v5110; shift_adder #(21, 14, 1, 1, 23, 8, 0) op_5110 (v2751[20:0], v3590[13:0], v5110[22:0]); // 4.0
    wire [24:0] v5111; shift_adder #(25, 14, 1, 1, 25, 9, 0) op_5111 (v3591[24:0], v3592[13:0], v5111[24:0]); // 4.0
    wire [26:0] v5112; shift_adder #(11, 27, 1, 1, 27, 0, 1) op_5112 (v237[10:0], v3593[26:0], v5112[26:0]); // 4.0
    wire [14:0] v5113; shift_adder #(13, 12, 1, 1, 15, 2, 0) op_5113 (v3594[12:0], v3595[11:0], v5113[14:0]); // 4.0
    wire [25:0] v5114; shift_adder #(16, 25, 1, 1, 26, -9, 0) op_5114 (v3596[15:0], v3597[24:0], v5114[25:0]); // 4.0
    wire [16:0] v5115; shift_adder #(15, 14, 1, 1, 17, 3, 0) op_5115 (v3598[14:0], v3599[13:0], v5115[16:0]); // 4.0
    wire [20:0] v5116; shift_adder #(18, 19, 1, 1, 21, -2, 0) op_5116 (v3600[17:0], v3404[18:0], v5116[20:0]); // 4.0
    wire [17:0] v5117; shift_adder #(17, 16, 1, 1, 18, 0, 0) op_5117 (v3601[16:0], v3602[15:0], v5117[17:0]); // 4.0
    wire [16:0] v5118; shift_adder #(15, 14, 1, 1, 17, 3, 0) op_5118 (v3603[14:0], v3604[13:0], v5118[16:0]); // 4.0
    wire [33:0] v5119; shift_adder #(32, 34, 1, 1, 34, -1, 0) op_5119 (v3311[31:0], v3606[33:0], v5119[33:0]); // 4.0
    wire [28:0] v5120; shift_adder #(22, 29, 1, 1, 29, -6, 0) op_5120 (v3607[21:0], v2568[28:0], v5120[28:0]); // 4.0
    wire [23:0] v5121; shift_adder #(19, 23, 1, 1, 24, -3, 0) op_5121 (v2668[18:0], v3608[22:0], v5121[23:0]); // 4.0
    wire [36:0] v5122; shift_adder #(14, 13, 1, 1, 37, 24, 1) op_5122 (v3609[13:0], v1518[12:0], v5122[36:0]); // 4.0
    wire [40:0] v5123; shift_adder #(40, 13, 1, 1, 41, 27, 0) op_5123 (v3610[39:0], v3611[12:0], v5123[40:0]); // 4.0
    wire [37:0] v5124; shift_adder #(15, 37, 1, 1, 38, -23, 0) op_5124 (v3612[14:0], v3613[36:0], v5124[37:0]); // 4.0
    wire [19:0] v5125; shift_adder #(18, 19, 1, 1, 20, -2, 0) op_5125 (v3614[17:0], v3615[18:0], v5125[19:0]); // 4.0
    wire [16:0] v5126; shift_adder #(17, 15, 1, 1, 17, 0, 0) op_5126 (v3181[16:0], v3616[14:0], v5126[16:0]); // 4.0
    wire [15:0] v5127; shift_adder #(14, 16, 1, 1, 16, -1, 0) op_5127 (v3617[13:0], v3618[15:0], v5127[15:0]); // 4.0
    wire [24:0] v5128; shift_adder #(8, 19, 1, 1, 25, -16, 1) op_5128 (v117[7:0], v3619[18:0], v5128[24:0]); // 4.0
    wire [22:0] v5129; shift_adder #(23, 16, 1, 1, 23, 6, 0) op_5129 (v3620[22:0], v3621[15:0], v5129[22:0]); // 4.0
    wire [28:0] v5130; shift_adder #(23, 27, 1, 1, 29, -6, 0) op_5130 (v3339[22:0], v3622[26:0], v5130[28:0]); // 4.0
    wire [24:0] v5131; shift_adder #(25, 23, 1, 1, 25, 0, 0) op_5131 (v3623[24:0], v3176[22:0], v5131[24:0]); // 4.0
    wire [24:0] v5132; shift_adder #(11, 23, 1, 1, 25, 2, 1) op_5132 (v201[10:0], v3624[22:0], v5132[24:0]); // 4.0
    wire [27:0] v5133; shift_adder #(18, 27, 1, 1, 28, -9, 0) op_5133 (v3625[17:0], v3317[26:0], v5133[27:0]); // 4.0
    wire [25:0] v5134; shift_adder #(26, 24, 1, 1, 26, 0, 0) op_5134 (v3626[25:0], v2899[23:0], v5134[25:0]); // 4.0
    wire [18:0] v5135; shift_adder #(17, 18, 1, 1, 19, -2, 0) op_5135 (v3627[16:0], v3628[17:0], v5135[18:0]); // 4.0
    wire [25:0] v5136; shift_adder #(17, 25, 1, 1, 26, -8, 0) op_5136 (v3629[16:0], v3630[24:0], v5136[25:0]); // 4.0
    wire [24:0] v5137; shift_adder #(25, 20, 1, 1, 25, 4, 0) op_5137 (v3457[24:0], v3554[19:0], v5137[24:0]); // 4.0
    wire [24:0] v5138; shift_adder #(18, 24, 1, 1, 25, -6, 0) op_5138 (v3631[17:0], v3632[23:0], v5138[24:0]); // 4.0
    wire [22:0] v5139; shift_adder #(21, 21, 1, 1, 23, -2, 0) op_5139 (v3633[20:0], v3634[20:0], v5139[22:0]); // 4.0
    wire [22:0] v5140; shift_adder #(18, 20, 1, 1, 23, -5, 0) op_5140 (v3635[17:0], v3292[19:0], v5140[22:0]); // 4.0
    wire [16:0] v5141; shift_adder #(16, 15, 1, 1, 17, 0, 0) op_5141 (v3636[15:0], v2704[14:0], v5141[16:0]); // 4.0
    wire [21:0] v5142; shift_adder #(18, 20, 1, 1, 22, -4, 0) op_5142 (v3637[17:0], v3237[19:0], v5142[21:0]); // 4.0
    wire [18:0] v5143; shift_adder #(12, 18, 1, 1, 19, -6, 1) op_5143 (v280[11:0], v3406[17:0], v5143[18:0]); // 4.0
    wire [21:0] v5144; shift_adder #(12, 22, 1, 1, 22, -9, 0) op_5144 (v3100[11:0], v3638[21:0], v5144[21:0]); // 4.0
    wire [21:0] v5145; shift_adder #(20, 20, 1, 1, 22, 1, 0) op_5145 (v3639[19:0], v3640[19:0], v5145[21:0]); // 4.0
    wire [22:0] v5146; shift_adder #(15, 23, 1, 1, 23, -7, 0) op_5146 (v3641[14:0], v3642[22:0], v5146[22:0]); // 4.0
    wire [21:0] v5147; shift_adder #(22, 13, 1, 1, 22, 7, 0) op_5147 (v2822[21:0], v3643[12:0], v5147[21:0]); // 4.0
    wire [29:0] v5148; shift_adder #(30, 25, 1, 1, 30, 4, 0) op_5148 (v3644[29:0], v3249[24:0], v5148[29:0]); // 4.0
    wire [25:0] v5149; shift_adder #(26, 19, 1, 1, 26, 6, 0) op_5149 (v3447[25:0], v3645[18:0], v5149[25:0]); // 4.0
    wire [21:0] v5150; shift_adder #(14, 20, 1, 1, 22, -7, 0) op_5150 (v3646[13:0], v2550[19:0], v5150[21:0]); // 4.0
    wire [18:0] v5151; shift_adder #(13, 18, 1, 1, 19, -5, 0) op_5151 (v3157[12:0], v3647[17:0], v5151[18:0]); // 4.0
    wire [28:0] v5152; shift_adder #(16, 28, 1, 1, 29, -12, 0) op_5152 (v3438[15:0], v3648[27:0], v5152[28:0]); // 4.0
    wire [34:0] v5153; shift_adder #(34, 13, 1, 1, 35, 21, 0) op_5153 (v3649[33:0], v3650[12:0], v5153[34:0]); // 4.0
    wire [18:0] v5154; shift_adder #(18, 16, 1, 1, 19, 2, 0) op_5154 (v3651[17:0], v3652[15:0], v5154[18:0]); // 4.0
    wire [24:0] v5155; shift_adder #(24, 14, 1, 1, 25, 9, 0) op_5155 (v3653[23:0], v3654[13:0], v5155[24:0]); // 4.0
    wire [15:0] v5156; shift_adder #(16, 13, 1, 1, 16, 2, 0) op_5156 (v3655[15:0], v2745[12:0], v5156[15:0]); // 4.0
    wire [30:0] v5157; shift_adder #(31, 17, 1, 1, 31, 11, 0) op_5157 (v3656[30:0], v3657[16:0], v5157[30:0]); // 4.0
    wire [33:0] v5158; shift_adder #(33, 19, 1, 1, 34, 14, 0) op_5158 (v3658[32:0], v3659[18:0], v5158[33:0]); // 4.0
    wire [19:0] v5159; shift_adder #(14, 20, 1, 1, 20, -5, 0) op_5159 (v3660[13:0], v3661[19:0], v5159[19:0]); // 4.0
    wire [14:0] v5160; shift_adder #(14, 14, 1, 1, 15, 0, 0) op_5160 (v3662[13:0], v3663[13:0], v5160[14:0]); // 4.0
    wire [16:0] v5161; shift_adder #(14, 14, 1, 1, 17, -2, 0) op_5161 (v2638[13:0], v3664[13:0], v5161[16:0]); // 4.0
    wire [19:0] v5162; shift_adder #(10, 20, 1, 1, 20, -4, 0) op_5162 (v446[9:0], v3665[19:0], v5162[19:0]); // 4.0
    wire [17:0] v5163; shift_adder #(15, 15, 1, 1, 18, -3, 0) op_5163 (v3666[14:0], v3186[14:0], v5163[17:0]); // 4.0
    wire [19:0] v5164; shift_adder #(16, 16, 1, 1, 20, -3, 0) op_5164 (v3667[15:0], v3668[15:0], v5164[19:0]); // 4.0
    wire [16:0] v5165; shift_adder #(16, 14, 1, 1, 17, 1, 0) op_5165 (v3038[15:0], v2907[13:0], v5165[16:0]); // 4.0
    wire [17:0] v5166; shift_adder #(17, 15, 1, 1, 18, 1, 0) op_5166 (v3569[16:0], v3669[14:0], v5166[17:0]); // 4.0
    wire [26:0] v5167; shift_adder #(11, 27, 1, 1, 27, -2, 1) op_5167 (v219[10:0], v3474[26:0], v5167[26:0]); // 4.0
    wire [25:0] v5168; shift_adder #(25, 18, 1, 1, 26, 8, 0) op_5168 (v3670[24:0], v3671[17:0], v5168[25:0]); // 4.0
    wire [26:0] v5169; shift_adder #(25, 27, 1, 1, 27, -1, 0) op_5169 (v3672[24:0], v3673[26:0], v5169[26:0]); // 4.0
    wire [19:0] v5170; shift_adder #(18, 18, 1, 1, 20, -2, 0) op_5170 (v3674[17:0], v2554[17:0], v5170[19:0]); // 4.0
    wire [20:0] v5171; shift_adder #(17, 21, 1, 1, 21, -3, 0) op_5171 (v3675[16:0], v3566[20:0], v5171[20:0]); // 4.0
    wire [24:0] v5172; shift_adder #(16, 23, 1, 1, 25, -9, 0) op_5172 (v2949[15:0], v3676[22:0], v5172[24:0]); // 4.0
    wire [25:0] v5173; shift_adder #(24, 18, 1, 1, 26, 7, 0) op_5173 (v3677[23:0], v3678[17:0], v5173[25:0]); // 4.0
    wire [25:0] v5174; shift_adder #(16, 25, 1, 1, 26, -9, 0) op_5174 (v3679[15:0], v3680[24:0], v5174[25:0]); // 4.0
    wire [30:0] v5175; shift_adder #(16, 30, 1, 1, 31, -11, 0) op_5175 (v3681[15:0], v3682[29:0], v5175[30:0]); // 4.0
    wire [30:0] v5176; shift_adder #(30, 31, 1, 1, 31, 0, 0) op_5176 (v3683[29:0], v3684[30:0], v5176[30:0]); // 4.0
    wire [21:0] v5177; shift_adder #(14, 21, 1, 1, 22, -7, 0) op_5177 (v3685[13:0], v3686[20:0], v5177[21:0]); // 4.0
    wire [26:0] v5178; shift_adder #(16, 16, 1, 1, 27, -11, 0) op_5178 (v3602[15:0], v3687[15:0], v5178[26:0]); // 4.0
    wire [32:0] v5179; shift_adder #(31, 20, 1, 1, 33, 12, 0) op_5179 (v2539[30:0], v3688[19:0], v5179[32:0]); // 4.0
    wire [17:0] v5180; shift_adder #(16, 17, 1, 1, 18, 0, 0) op_5180 (v3689[15:0], v3690[16:0], v5180[17:0]); // 4.0
    wire [18:0] v5181; shift_adder #(15, 19, 1, 1, 19, -1, 0) op_5181 (v3691[14:0], v3692[18:0], v5181[18:0]); // 4.0
    wire [14:0] v5182; shift_adder #(14, 13, 1, 1, 15, 0, 0) op_5182 (v3049[13:0], v3693[12:0], v5182[14:0]); // 4.0
    wire [33:0] v5183; shift_adder #(12, 13, 1, 1, 34, 21, 1) op_5183 (v2733[11:0], v2018[12:0], v5183[33:0]); // 4.0
    wire [14:0] v5184; shift_adder #(13, 13, 1, 1, 15, 1, 0) op_5184 (v2860[12:0], v3694[12:0], v5184[14:0]); // 4.0
    wire [17:0] v5185; shift_adder #(17, 15, 1, 1, 18, 2, 0) op_5185 (v3695[16:0], v3696[14:0], v5185[17:0]); // 4.0
    wire [25:0] v5186; shift_adder #(21, 25, 1, 1, 26, -4, 0) op_5186 (v3147[20:0], v3697[24:0], v5186[25:0]); // 4.0
    wire [23:0] v5187; shift_adder #(23, 19, 1, 1, 24, 4, 0) op_5187 (v3698[22:0], v3699[18:0], v5187[23:0]); // 4.0
    wire [22:0] v5188; shift_adder #(21, 22, 1, 1, 23, 1, 0) op_5188 (v3109[20:0], v3700[21:0], v5188[22:0]); // 4.0
    wire [15:0] v5189; shift_adder #(13, 16, 1, 1, 16, -1, 0) op_5189 (v3701[12:0], v3702[15:0], v5189[15:0]); // 4.0
    wire [26:0] v5190; shift_adder #(26, 22, 1, 1, 27, 5, 0) op_5190 (v3703[25:0], v2605[21:0], v5190[26:0]); // 4.0
    wire [27:0] v5191; shift_adder #(27, 18, 1, 1, 28, 10, 0) op_5191 (v3704[26:0], v3705[17:0], v5191[27:0]); // 4.0
    wire [18:0] v5192; shift_adder #(18, 16, 1, 1, 19, 2, 0) op_5192 (v2597[17:0], v3706[15:0], v5192[18:0]); // 4.0
    wire [26:0] v5193; shift_adder #(26, 17, 1, 1, 27, 9, 0) op_5193 (v3707[25:0], v3179[16:0], v5193[26:0]); // 4.0
    wire [22:0] v5194; shift_adder #(23, 15, 1, 1, 23, 7, 0) op_5194 (v3708[22:0], v2758[14:0], v5194[22:0]); // 4.0
    wire [21:0] v5195; shift_adder #(19, 21, 1, 1, 22, -2, 0) op_5195 (v3402[18:0], v3390[20:0], v5195[21:0]); // 4.0
    wire [33:0] v5196; shift_adder #(34, 29, 1, 1, 34, 3, 0) op_5196 (v3709[33:0], v3710[28:0], v5196[33:0]); // 4.0
    wire [13:0] v5197; shift_adder #(11, 14, 1, 1, 14, 0, 0) op_5197 (v144[10:0], v3711[13:0], v5197[13:0]); // 4.0
    wire [24:0] v5198; shift_adder #(24, 17, 1, 1, 25, 7, 0) op_5198 (v3712[23:0], v3713[16:0], v5198[24:0]); // 4.0
    wire [26:0] v5199; shift_adder #(21, 24, 1, 1, 27, -6, 0) op_5199 (v2767[20:0], v3714[23:0], v5199[26:0]); // 4.0
    wire [26:0] v5200; shift_adder #(15, 27, 1, 1, 27, -10, 1) op_5200 (v1473[14:0], v3715[26:0], v5200[26:0]); // 4.0
    wire [18:0] v5201; shift_adder #(15, 16, 1, 1, 19, 3, 0) op_5201 (v3716[14:0], v3717[15:0], v5201[18:0]); // 4.0
    wire [15:0] v5202; shift_adder #(14, 14, 1, 1, 16, 1, 0) op_5202 (v3662[13:0], v2574[13:0], v5202[15:0]); // 4.0
    wire [18:0] v5203; shift_adder #(18, 18, 1, 1, 19, 1, 0) op_5203 (v3718[17:0], v3719[17:0], v5203[18:0]); // 4.0
    wire [20:0] v5204; shift_adder #(11, 21, 1, 1, 21, -3, 1) op_5204 (v223[10:0], v3720[20:0], v5204[20:0]); // 4.0
    wire [22:0] v5205; shift_adder #(16, 22, 1, 1, 23, -6, 0) op_5205 (v3721[15:0], v3722[21:0], v5205[22:0]); // 4.0
    wire [34:0] v5206; shift_adder #(35, 17, 1, 1, 35, 17, 0) op_5206 (v3723[34:0], v3724[16:0], v5206[34:0]); // 4.0
    wire [27:0] v5207; shift_adder #(14, 28, 1, 1, 28, 0, 1) op_5207 (v499[13:0], v3725[27:0], v5207[27:0]); // 4.0
    wire [24:0] v5208; shift_adder #(24, 14, 1, 1, 25, 10, 0) op_5208 (v3726[23:0], v3727[13:0], v5208[24:0]); // 4.0
    wire [17:0] v5209; shift_adder #(15, 17, 1, 1, 18, -3, 0) op_5209 (v3345[14:0], v3519[16:0], v5209[17:0]); // 4.0
    wire [17:0] v5210; shift_adder #(15, 17, 1, 1, 18, -2, 0) op_5210 (v3728[14:0], v3729[16:0], v5210[17:0]); // 4.0
    wire [23:0] v5211; shift_adder #(16, 23, 1, 1, 24, -7, 0) op_5211 (v2564[15:0], v3320[22:0], v5211[23:0]); // 4.0
    wire [25:0] v5212; shift_adder #(25, 21, 1, 1, 26, 2, 0) op_5212 (v3730[24:0], v3731[20:0], v5212[25:0]); // 4.0
    wire [20:0] v5213; shift_adder #(18, 19, 1, 1, 21, -3, 0) op_5213 (v2640[17:0], v3732[18:0], v5213[20:0]); // 4.0
    wire [19:0] v5214; shift_adder #(17, 20, 1, 1, 20, -1, 0) op_5214 (v3733[16:0], v3734[19:0], v5214[19:0]); // 4.0
    wire [25:0] v5215; shift_adder #(13, 18, 1, 1, 26, -13, 0) op_5215 (v578[12:0], v3097[17:0], v5215[25:0]); // 4.0
    wire [37:0] v5216; shift_adder #(37, 31, 1, 1, 38, 5, 0) op_5216 (v3735[36:0], v3736[30:0], v5216[37:0]); // 4.0
    wire [23:0] v5217; shift_adder #(23, 21, 1, 1, 24, 3, 0) op_5217 (v3737[22:0], v3403[20:0], v5217[23:0]); // 4.0
    wire [24:0] v5218; shift_adder #(15, 24, 1, 1, 25, -9, 0) op_5218 (v3738[14:0], v3739[23:0], v5218[24:0]); // 4.0
    wire [33:0] v5219; shift_adder #(33, 31, 1, 1, 34, 3, 0) op_5219 (v3740[32:0], v3003[30:0], v5219[33:0]); // 4.0
    wire [30:0] v5220; shift_adder #(30, 16, 1, 1, 31, 15, 0) op_5220 (v3741[29:0], v3742[15:0], v5220[30:0]); // 4.0
    wire [37:0] v5221; shift_adder #(20, 38, 1, 1, 38, -16, 0) op_5221 (v3743[19:0], v3744[37:0], v5221[37:0]); // 4.0
    wire [16:0] v5222; shift_adder #(14, 16, 1, 1, 17, -2, 0) op_5222 (v3745[13:0], v3746[15:0], v5222[16:0]); // 4.0
    wire [16:0] v5223; shift_adder #(17, 15, 1, 1, 17, 1, 0) op_5223 (v3747[16:0], v3748[14:0], v5223[16:0]); // 4.0
    wire [15:0] v5224; shift_adder #(14, 14, 1, 1, 16, 1, 0) op_5224 (v3749[13:0], v3750[13:0], v5224[15:0]); // 4.0
    wire [20:0] v5225; shift_adder #(13, 21, 1, 1, 21, -7, 1) op_5225 (v932[12:0], v3751[20:0], v5225[20:0]); // 4.0
    wire [19:0] v5226; shift_adder #(18, 15, 1, 1, 20, 4, 0) op_5226 (v3752[17:0], v2894[14:0], v5226[19:0]); // 4.0
    wire [20:0] v5227; shift_adder #(19, 19, 1, 1, 21, -1, 0) op_5227 (v3753[18:0], v3117[18:0], v5227[20:0]); // 4.0
    wire [20:0] v5228; shift_adder #(18, 20, 1, 1, 21, -2, 0) op_5228 (v3754[17:0], v3755[19:0], v5228[20:0]); // 4.0
    wire [18:0] v5229; shift_adder #(16, 18, 1, 1, 19, -3, 1) op_5229 (v2685[15:0], v562[17:0], v5229[18:0]); // 4.0
    wire [22:0] v5230; shift_adder #(16, 22, 1, 1, 23, -4, 0) op_5230 (v3756[15:0], v3757[21:0], v5230[22:0]); // 4.0
    wire [22:0] v5231; shift_adder #(21, 22, 1, 1, 23, -1, 0) op_5231 (v3758[20:0], v3759[21:0], v5231[22:0]); // 4.0
    wire [23:0] v5232; shift_adder #(17, 23, 1, 1, 24, -6, 0) op_5232 (v3760[16:0], v3761[22:0], v5232[23:0]); // 4.0
    wire [21:0] v5233; shift_adder #(21, 15, 1, 1, 22, 6, 0) op_5233 (v3552[20:0], v3762[14:0], v5233[21:0]); // 4.0
    wire [25:0] v5234; shift_adder #(13, 26, 1, 1, 26, -12, 0) op_5234 (v3763[12:0], v3506[25:0], v5234[25:0]); // 4.0
    wire [25:0] v5235; shift_adder #(25, 20, 1, 1, 26, 4, 0) op_5235 (v3350[24:0], v3764[19:0], v5235[25:0]); // 4.0
    wire [24:0] v5236; shift_adder #(16, 24, 1, 1, 25, -7, 0) op_5236 (v3765[15:0], v3766[23:0], v5236[24:0]); // 4.0
    wire [29:0] v5237; shift_adder #(29, 14, 1, 1, 30, 15, 0) op_5237 (v3767[28:0], v3768[13:0], v5237[29:0]); // 4.0
    wire [27:0] v5238; shift_adder #(15, 27, 1, 1, 28, -11, 0) op_5238 (v2625[14:0], v3769[26:0], v5238[27:0]); // 4.0
    wire [28:0] v5239; shift_adder #(15, 28, 1, 1, 29, -13, 0) op_5239 (v3105[14:0], v2525[27:0], v5239[28:0]); // 4.0
    wire [25:0] v5240; shift_adder #(25, 17, 1, 1, 26, 9, 0) op_5240 (v3770[24:0], v3771[16:0], v5240[25:0]); // 4.0
    wire [17:0] v5241; shift_adder #(14, 18, 1, 1, 18, 0, 0) op_5241 (v3772[13:0], v2650[17:0], v5241[17:0]); // 4.0
    wire [15:0] v5242; shift_adder #(15, 14, 1, 1, 16, 1, 0) op_5242 (v3773[14:0], v3106[13:0], v5242[15:0]); // 4.0
    wire [20:0] v5243; shift_adder #(20, 17, 1, 1, 21, 3, 0) op_5243 (v3774[19:0], v3775[16:0], v5243[20:0]); // 4.0
    wire [22:0] v5244; shift_adder #(21, 19, 1, 1, 23, 4, 0) op_5244 (v3776[20:0], v3220[18:0], v5244[22:0]); // 4.0
    wire [20:0] v5245; shift_adder #(20, 15, 1, 1, 21, 4, 0) op_5245 (v3777[19:0], v3778[14:0], v5245[20:0]); // 4.0
    wire [20:0] v5246; shift_adder #(21, 15, 1, 1, 21, 2, 0) op_5246 (v3779[20:0], v2794[14:0], v5246[20:0]); // 4.0
    wire [14:0] v5247; shift_adder #(14, 13, 1, 1, 15, -1, 0) op_5247 (v3780[13:0], v3781[12:0], v5247[14:0]); // 4.0
    wire [31:0] v5248; shift_adder #(32, 14, 1, 1, 32, 17, 0) op_5248 (v3782[31:0], v3061[13:0], v5248[31:0]); // 4.0
    wire [29:0] v5249; shift_adder #(29, 23, 1, 1, 30, 6, 0) op_5249 (v3783[28:0], v3784[22:0], v5249[29:0]); // 4.0
    wire [35:0] v5250; shift_adder #(20, 14, 1, 1, 36, -16, 1) op_5250 (v3785[19:0], v3786[13:0], v5250[35:0]); // 4.0
    wire [35:0] v5251; shift_adder #(35, 35, 1, 1, 36, 0, 0) op_5251 (v3787[34:0], v3788[34:0], v5251[35:0]); // 4.0
    wire [24:0] v5252; shift_adder #(24, 21, 1, 1, 25, 3, 0) op_5252 (v2553[23:0], v3789[20:0], v5252[24:0]); // 4.0
    wire [37:0] v5253; shift_adder #(15, 36, 1, 1, 38, -22, 0) op_5253 (v3790[14:0], v3791[35:0], v5253[37:0]); // 4.0
    wire [33:0] v5254; shift_adder #(33, 25, 1, 1, 34, 9, 0) op_5254 (v3299[32:0], v3570[24:0], v5254[33:0]); // 4.0
    wire [23:0] v5255; shift_adder #(16, 22, 1, 1, 24, -7, 0) op_5255 (v3792[15:0], v2621[21:0], v5255[23:0]); // 4.0
    wire [29:0] v5256; shift_adder #(29, 17, 1, 1, 30, 11, 0) op_5256 (v3793[28:0], v3794[16:0], v5256[29:0]); // 4.0
    wire [26:0] v5257; shift_adder #(11, 23, 1, 1, 27, -16, 0) op_5257 (v155[10:0], v3795[22:0], v5257[26:0]); // 4.0
    wire [16:0] v5258; shift_adder #(16, 16, 1, 1, 17, 0, 0) op_5258 (v3796[15:0], v3797[15:0], v5258[16:0]); // 4.0
    wire [27:0] v5259; shift_adder #(27, 20, 1, 1, 28, 7, 0) op_5259 (v3503[26:0], v3798[19:0], v5259[27:0]); // 4.0
    wire [16:0] v5260; shift_adder #(16, 16, 1, 1, 17, 0, 0) op_5260 (v3799[15:0], v3800[15:0], v5260[16:0]); // 4.0
    wire [25:0] v5261; shift_adder #(26, 20, 1, 1, 26, 2, 0) op_5261 (v3801[25:0], v3802[19:0], v5261[25:0]); // 4.0
    wire [29:0] v5262; shift_adder #(29, 26, 1, 1, 30, 3, 0) op_5262 (v3185[28:0], v3020[25:0], v5262[29:0]); // 4.0
    wire [26:0] v5263; shift_adder #(13, 27, 1, 1, 27, -13, 0) op_5263 (v3803[12:0], v3804[26:0], v5263[26:0]); // 4.0
    wire [28:0] v5264; shift_adder #(25, 28, 1, 1, 29, -3, 0) op_5264 (v3805[24:0], v3806[27:0], v5264[28:0]); // 4.0
    wire [24:0] v5265; shift_adder #(24, 22, 1, 1, 25, 3, 0) op_5265 (v3807[23:0], v3808[21:0], v5265[24:0]); // 4.0
    wire [17:0] v5266; shift_adder #(16, 16, 1, 1, 18, 2, 0) op_5266 (v3809[15:0], v3810[15:0], v5266[17:0]); // 4.0
    wire [22:0] v5267; shift_adder #(13, 23, 1, 1, 23, -2, 1) op_5267 (v932[12:0], v3811[22:0], v5267[22:0]); // 4.0
    wire [24:0] v5268; shift_adder #(24, 22, 1, 1, 25, 1, 0) op_5268 (v3812[23:0], v3813[21:0], v5268[24:0]); // 4.0
    wire [22:0] v5269; shift_adder #(16, 23, 1, 1, 23, -5, 0) op_5269 (v3814[15:0], v3815[22:0], v5269[22:0]); // 4.0
    wire [17:0] v5270; shift_adder #(16, 14, 1, 1, 18, 3, 0) op_5270 (v3816[15:0], v2818[13:0], v5270[17:0]); // 4.0
    wire [19:0] v5271; shift_adder #(18, 17, 1, 1, 20, 3, 0) op_5271 (v3817[17:0], v3818[16:0], v5271[19:0]); // 4.0
    wire [21:0] v5272; shift_adder #(14, 22, 1, 1, 22, -6, 0) op_5272 (v3149[13:0], v3819[21:0], v5272[21:0]); // 4.0
    wire [24:0] v5273; shift_adder #(22, 24, 1, 1, 25, 1, 0) op_5273 (v2924[21:0], v3364[23:0], v5273[24:0]); // 4.0
    wire [20:0] v5274; shift_adder #(16, 20, 1, 1, 21, -4, 0) op_5274 (v3820[15:0], v3163[19:0], v5274[20:0]); // 4.0
    wire [24:0] v5275; shift_adder #(24, 22, 1, 1, 25, 2, 0) op_5275 (v3821[23:0], v3822[21:0], v5275[24:0]); // 4.0
    wire [25:0] v5276; shift_adder #(12, 19, 1, 1, 26, -14, 1) op_5276 (v2116[11:0], v3823[18:0], v5276[25:0]); // 4.0
    wire [24:0] v5277; shift_adder #(24, 19, 1, 1, 25, 5, 0) op_5277 (v3824[23:0], v3825[18:0], v5277[24:0]); // 4.0
    wire [25:0] v5278; shift_adder #(18, 25, 1, 1, 26, -6, 0) op_5278 (v2749[17:0], v3134[24:0], v5278[25:0]); // 4.0
    wire [26:0] v5279; shift_adder #(20, 26, 1, 1, 27, -6, 0) op_5279 (v3826[19:0], v2756[25:0], v5279[26:0]); // 4.0
    wire [25:0] v5280; shift_adder #(23, 19, 1, 1, 26, 6, 0) op_5280 (v3827[22:0], v3828[18:0], v5280[25:0]); // 4.0
    wire [31:0] v5281; shift_adder #(30, 28, 1, 1, 32, 3, 0) op_5281 (v3683[29:0], v3564[27:0], v5281[31:0]); // 4.0
    wire [23:0] v5282; shift_adder #(22, 23, 1, 1, 24, -1, 0) op_5282 (v3829[21:0], v3737[22:0], v5282[23:0]); // 4.0
    wire [30:0] v5283; shift_adder #(30, 16, 1, 1, 31, 13, 0) op_5283 (v3830[29:0], v3831[15:0], v5283[30:0]); // 4.0
    wire [36:0] v5284; shift_adder #(37, 15, 1, 1, 37, 21, 0) op_5284 (v3832[36:0], v3833[14:0], v5284[36:0]); // 4.0
    wire [15:0] v5285; shift_adder #(14, 15, 1, 1, 16, -1, 0) op_5285 (v3834[13:0], v3835[14:0], v5285[15:0]); // 4.0
    wire [38:0] v5286; shift_adder #(33, 38, 1, 1, 39, -4, 0) op_5286 (v3836[32:0], v3837[37:0], v5286[38:0]); // 4.0
    wire [38:0] v5287; shift_adder #(16, 15, 1, 1, 39, 24, 1) op_5287 (v3838[15:0], v945[14:0], v5287[38:0]); // 4.0
    wire [23:0] v5288; shift_adder #(15, 21, 1, 1, 24, -8, 0) op_5288 (v3839[14:0], v3840[20:0], v5288[23:0]); // 4.0
    wire [22:0] v5289; shift_adder #(17, 21, 1, 1, 23, -5, 0) op_5289 (v3841[16:0], v3842[20:0], v5289[22:0]); // 4.0
    wire [16:0] v5290; shift_adder #(16, 15, 1, 1, 17, -1, 0) op_5290 (v2952[15:0], v3843[14:0], v5290[16:0]); // 4.0
    wire [16:0] v5291; shift_adder #(15, 15, 1, 1, 17, -1, 0) op_5291 (v3844[14:0], v3845[14:0], v5291[16:0]); // 4.0
    wire [18:0] v5292; shift_adder #(15, 16, 1, 1, 19, 3, 0) op_5292 (v3846[14:0], v3847[15:0], v5292[18:0]); // 4.0
    wire [18:0] v5293; shift_adder #(15, 18, 1, 1, 19, -2, 0) op_5293 (v3848[14:0], v3849[17:0], v5293[18:0]); // 4.0
    wire [26:0] v5294; shift_adder #(26, 23, 1, 1, 27, 3, 0) op_5294 (v3850[25:0], v3851[22:0], v5294[26:0]); // 4.0
    wire [32:0] v5295; shift_adder #(32, 16, 1, 1, 33, 16, 0) op_5295 (v3560[31:0], v3852[15:0], v5295[32:0]); // 4.0
    wire [22:0] v5296; shift_adder #(14, 22, 1, 1, 23, -8, 0) op_5296 (v3853[13:0], v3530[21:0], v5296[22:0]); // 4.0
    wire [26:0] v5297; shift_adder #(19, 26, 1, 1, 27, -7, 0) op_5297 (v3854[18:0], v3855[25:0], v5297[26:0]); // 4.0
    wire [19:0] v5298; shift_adder #(13, 19, 1, 1, 20, -6, 0) op_5298 (v3701[12:0], v3856[18:0], v5298[19:0]); // 4.0
    wire [27:0] v5299; shift_adder #(27, 15, 1, 1, 28, 12, 0) op_5299 (v3804[26:0], v3857[14:0], v5299[27:0]); // 4.0
    wire [23:0] v5300; shift_adder #(23, 14, 1, 1, 24, 9, 0) op_5300 (v3327[22:0], v3858[13:0], v5300[23:0]); // 4.0
    wire [28:0] v5301; shift_adder #(27, 25, 1, 1, 29, 4, 0) op_5301 (v3077[26:0], v3229[24:0], v5301[28:0]); // 4.0
    wire [31:0] v5302; shift_adder #(32, 16, 1, 1, 32, 12, 0) op_5302 (v3859[31:0], v3860[15:0], v5302[31:0]); // 4.0
    wire [32:0] v5303; shift_adder #(33, 28, 1, 1, 33, 4, 0) op_5303 (v2930[32:0], v3559[27:0], v5303[32:0]); // 4.0
    wire [24:0] v5304; shift_adder #(16, 23, 1, 1, 25, -8, 0) op_5304 (v2916[15:0], v3861[22:0], v5304[24:0]); // 4.0
    wire [32:0] v5305; shift_adder #(33, 28, 1, 1, 33, 3, 0) op_5305 (v3862[32:0], v3863[27:0], v5305[32:0]); // 4.0
    wire [17:0] v5306; shift_adder #(15, 17, 1, 1, 18, -2, 0) op_5306 (v3864[14:0], v2801[16:0], v5306[17:0]); // 4.0
    wire [22:0] v5307; shift_adder #(22, 16, 1, 1, 23, 6, 0) op_5307 (v3516[21:0], v3865[15:0], v5307[22:0]); // 4.0
    wire [26:0] v5308; shift_adder #(26, 17, 1, 1, 27, 9, 0) op_5308 (v3866[25:0], v3867[16:0], v5308[26:0]); // 4.0
    wire [25:0] v5309; shift_adder #(26, 16, 1, 1, 26, 7, 0) op_5309 (v3868[25:0], v3869[15:0], v5309[25:0]); // 4.0
    wire [29:0] v5310; shift_adder #(30, 15, 1, 1, 30, 12, 0) op_5310 (v3870[29:0], v3871[14:0], v5310[29:0]); // 4.0
    wire [21:0] v5311; shift_adder #(17, 21, 1, 1, 22, -4, 0) op_5311 (v3872[16:0], v3873[20:0], v5311[21:0]); // 4.0
    wire [22:0] v5312; shift_adder #(18, 22, 1, 1, 23, -3, 0) op_5312 (v2764[17:0], v3874[21:0], v5312[22:0]); // 4.0
    wire [17:0] v5313; shift_adder #(17, 13, 1, 1, 18, 4, 0) op_5313 (v3875[16:0], v2528[12:0], v5313[17:0]); // 4.0
    wire [20:0] v5314; shift_adder #(15, 21, 1, 1, 21, -5, 0) op_5314 (v2865[14:0], v3876[20:0], v5314[20:0]); // 4.0
    wire [26:0] v5315; shift_adder #(14, 27, 1, 1, 27, -10, 0) op_5315 (v3654[13:0], v3877[26:0], v5315[26:0]); // 4.0
    wire [27:0] v5316; shift_adder #(25, 19, 1, 1, 28, 9, 0) op_5316 (v3878[24:0], v3879[18:0], v5316[27:0]); // 4.0
    wire [34:0] v5317; shift_adder #(29, 35, 1, 1, 35, -5, 0) op_5317 (v3880[28:0], v3881[34:0], v5317[34:0]); // 4.0
    wire [17:0] v5318; shift_adder #(14, 17, 1, 1, 18, 1, 0) op_5318 (v3882[13:0], v3883[16:0], v5318[17:0]); // 4.0
    wire [17:0] v5319; shift_adder #(16, 17, 1, 1, 18, 0, 0) op_5319 (v3884[15:0], v3885[16:0], v5319[17:0]); // 4.0
    wire [24:0] v5320; shift_adder #(23, 23, 1, 1, 25, -2, 0) op_5320 (v2771[22:0], v3123[22:0], v5320[24:0]); // 4.0
    wire [18:0] v5321; shift_adder #(17, 16, 1, 1, 19, 3, 0) op_5321 (v3886[16:0], v3887[15:0], v5321[18:0]); // 4.0
    wire [35:0] v5322; shift_adder #(13, 35, 1, 1, 36, -22, 0) op_5322 (v3888[12:0], v3723[34:0], v5322[35:0]); // 4.0
    wire [22:0] v5323; shift_adder #(20, 21, 1, 1, 23, -2, 0) op_5323 (v3023[19:0], v2716[20:0], v5323[22:0]); // 4.0
    wire [31:0] v5324; shift_adder #(31, 19, 1, 1, 32, 12, 0) op_5324 (v3890[30:0], v3891[18:0], v5324[31:0]); // 4.0
    wire [27:0] v5325; shift_adder #(27, 24, 1, 1, 28, 3, 0) op_5325 (v3892[26:0], v3893[23:0], v5325[27:0]); // 4.0
    wire [20:0] v5326; shift_adder #(20, 18, 1, 1, 21, 2, 0) op_5326 (v3894[19:0], v3164[17:0], v5326[20:0]); // 4.0
    wire [29:0] v5327; shift_adder #(29, 28, 1, 1, 30, 2, 0) op_5327 (v2824[28:0], v3563[27:0], v5327[29:0]); // 4.0
    wire [38:0] v5328; shift_adder #(17, 12, 1, 1, 39, 27, 1) op_5328 (v3895[16:0], v2077[11:0], v5328[38:0]); // 4.0
    wire [36:0] v5329; shift_adder #(35, 15, 1, 1, 37, -2, 1) op_5329 (v3896[34:0], v3897[14:0], v5329[36:0]); // 4.0
    wire [36:0] v5330; shift_adder #(35, 14, 1, 1, 37, 22, 0) op_5330 (v3898[34:0], v3899[13:0], v5330[36:0]); // 4.0
    wire [20:0] v5331; shift_adder #(20, 19, 1, 1, 21, -1, 0) op_5331 (v3576[19:0], v3900[18:0], v5331[20:0]); // 4.0
    wire [18:0] v5332; shift_adder #(17, 17, 1, 1, 19, -1, 0) op_5332 (v2920[16:0], v3901[16:0], v5332[18:0]); // 4.0
    wire [15:0] v5333; shift_adder #(15, 14, 1, 1, 16, 1, 0) op_5333 (v3902[14:0], v3903[13:0], v5333[15:0]); // 4.0
    wire [18:0] v5334; shift_adder #(18, 16, 1, 1, 19, 2, 0) op_5334 (v3904[17:0], v3312[15:0], v5334[18:0]); // 4.0
    wire [20:0] v5335; shift_adder #(20, 13, 1, 1, 21, 6, 0) op_5335 (v3905[19:0], v3906[12:0], v5335[20:0]); // 4.0
    wire [33:0] v5336; shift_adder #(34, 23, 1, 1, 34, 9, 0) op_5336 (v3907[33:0], v3908[22:0], v5336[33:0]); // 4.0
    wire [26:0] v5337; shift_adder #(27, 21, 1, 1, 27, 4, 0) op_5337 (v2620[26:0], v3909[20:0], v5337[26:0]); // 4.0
    wire [31:0] v5338; shift_adder #(22, 31, 1, 1, 32, -10, 0) op_5338 (v3526[21:0], v3910[30:0], v5338[31:0]); // 4.0
    wire [21:0] v5339; shift_adder #(21, 19, 1, 1, 22, -1, 0) op_5339 (v2648[20:0], v3911[18:0], v5339[21:0]); // 4.0
    wire [25:0] v5340; shift_adder #(26, 17, 1, 1, 26, 7, 0) op_5340 (v3912[25:0], v3913[16:0], v5340[25:0]); // 4.0
    wire [17:0] v5341; shift_adder #(15, 16, 1, 1, 18, -3, 0) op_5341 (v3914[14:0], v3915[15:0], v5341[17:0]); // 4.0
    wire [22:0] v5342; shift_adder #(12, 23, 1, 1, 23, -7, 1) op_5342 (v999[11:0], v3916[22:0], v5342[22:0]); // 4.0
    wire [18:0] v5343; shift_adder #(19, 16, 1, 1, 19, 2, 0) op_5343 (v3917[18:0], v3918[15:0], v5343[18:0]); // 4.0
    wire [17:0] v5344; shift_adder #(18, 16, 1, 1, 18, 1, 0) op_5344 (v3489[17:0], v3919[15:0], v5344[17:0]); // 4.0
    wire [21:0] v5345; shift_adder #(22, 16, 1, 1, 22, 4, 0) op_5345 (v3700[21:0], v3920[15:0], v5345[21:0]); // 4.0
    wire [21:0] v5346; shift_adder #(21, 14, 1, 1, 22, 6, 0) op_5346 (v2897[20:0], v3921[13:0], v5346[21:0]); // 4.0
    wire [16:0] v5347; shift_adder #(17, 14, 1, 1, 17, 1, 0) op_5347 (v3922[16:0], v3923[13:0], v5347[16:0]); // 4.0
    wire [20:0] v5348; shift_adder #(20, 15, 1, 1, 21, 6, 0) op_5348 (v3924[19:0], v3925[14:0], v5348[20:0]); // 4.0
    wire [18:0] v5349; shift_adder #(18, 15, 1, 1, 19, 4, 0) op_5349 (v3129[17:0], v3926[14:0], v5349[18:0]); // 4.0
    wire [19:0] v5350; shift_adder #(15, 19, 1, 1, 20, -3, 0) op_5350 (v3927[14:0], v3413[18:0], v5350[19:0]); // 4.0
    wire [24:0] v5351; shift_adder #(18, 24, 1, 1, 25, -6, 0) op_5351 (v3928[17:0], v3929[23:0], v5351[24:0]); // 4.0
    wire [29:0] v5352; shift_adder #(18, 29, 1, 1, 30, -10, 0) op_5352 (v3637[17:0], v3930[28:0], v5352[29:0]); // 4.0
    wire [22:0] v5353; shift_adder #(21, 22, 1, 1, 23, 0, 0) op_5353 (v3931[20:0], v3932[21:0], v5353[22:0]); // 4.0
    wire [20:0] v5354; shift_adder #(15, 20, 1, 1, 21, -4, 0) op_5354 (v2694[14:0], v3323[19:0], v5354[20:0]); // 4.0
    wire [17:0] v5355; shift_adder #(16, 16, 1, 1, 18, 1, 0) op_5355 (v3933[15:0], v3934[15:0], v5355[17:0]); // 4.0
    wire [25:0] v5356; shift_adder #(18, 26, 1, 1, 26, -4, 0) op_5356 (v3935[17:0], v3936[25:0], v5356[25:0]); // 4.0
    wire [21:0] v5357; shift_adder #(22, 16, 1, 1, 22, 5, 0) op_5357 (v2993[21:0], v3937[15:0], v5357[21:0]); // 4.0
    wire [30:0] v5358; shift_adder #(31, 15, 1, 1, 31, 15, 0) op_5358 (v3938[30:0], v3939[14:0], v5358[30:0]); // 4.0
    wire [14:0] v5359; shift_adder #(12, 15, 1, 1, 15, 0, 0) op_5359 (v3417[11:0], v3346[14:0], v5359[14:0]); // 4.0
    wire [18:0] v5360; shift_adder #(17, 14, 1, 1, 19, 4, 0) op_5360 (v3940[16:0], v3941[13:0], v5360[18:0]); // 4.0
    wire [35:0] v5361; shift_adder #(16, 35, 1, 1, 36, -20, 0) op_5361 (v3942[15:0], v3943[34:0], v5361[35:0]); // 4.0
    wire [39:0] v5362; shift_adder #(15, 38, 1, 1, 40, -24, 0) op_5362 (v3641[14:0], v3944[37:0], v5362[39:0]); // 4.0
    wire [22:0] v5363; shift_adder #(22, 18, 1, 1, 23, 4, 0) op_5363 (v3449[21:0], v3945[17:0], v5363[22:0]); // 4.0
    wire [36:0] v5364; shift_adder #(16, 36, 1, 1, 37, -20, 0) op_5364 (v3946[15:0], v3947[35:0], v5364[36:0]); // 4.0
    wire [13:0] v5365; shift_adder #(14, 13, 1, 1, 14, 0, 0) op_5365 (v3948[13:0], v2975[12:0], v5365[13:0]); // 4.0
    wire [25:0] v5366; shift_adder #(19, 24, 1, 1, 26, -6, 0) op_5366 (v3949[18:0], v3950[23:0], v5366[25:0]); // 4.0
    wire [16:0] v5367; shift_adder #(14, 16, 1, 1, 17, -2, 0) op_5367 (v3951[13:0], v3706[15:0], v5367[16:0]); // 4.0
    wire [19:0] v5368; shift_adder #(11, 20, 1, 1, 20, -6, 0) op_5368 (v323[10:0], v3952[19:0], v5368[19:0]); // 4.0
    wire [20:0] v5369; shift_adder #(19, 20, 1, 1, 21, -2, 0) op_5369 (v3953[18:0], v3954[19:0], v5369[20:0]); // 4.0
    wire [17:0] v5370; shift_adder #(15, 16, 1, 1, 18, -3, 0) op_5370 (v3955[14:0], v3495[15:0], v5370[17:0]); // 4.0
    wire [17:0] v5371; shift_adder #(15, 16, 1, 1, 18, -2, 0) op_5371 (v3956[14:0], v3546[15:0], v5371[17:0]); // 4.0
    wire [21:0] v5372; shift_adder #(20, 16, 1, 1, 22, 5, 0) op_5372 (v3410[19:0], v3957[15:0], v5372[21:0]); // 4.0
    wire [28:0] v5373; shift_adder #(27, 27, 1, 1, 29, -1, 0) op_5373 (v3958[26:0], v3959[26:0], v5373[28:0]); // 4.0
    wire [15:0] v5374; shift_adder #(15, 15, 1, 1, 16, 0, 0) op_5374 (v2747[14:0], v3960[14:0], v5374[15:0]); // 4.0
    wire [22:0] v5375; shift_adder #(22, 20, 1, 1, 23, 2, 0) op_5375 (v3961[21:0], v3962[19:0], v5375[22:0]); // 4.0
    wire [17:0] v5376; shift_adder #(17, 16, 1, 1, 18, 1, 0) op_5376 (v3152[16:0], v3963[15:0], v5376[17:0]); // 4.0
    wire [16:0] v5377; shift_adder #(13, 16, 1, 1, 17, -2, 0) op_5377 (v3964[12:0], v3965[15:0], v5377[16:0]); // 4.0
    wire [28:0] v5378; shift_adder #(28, 22, 1, 1, 29, 7, 0) op_5378 (v3415[27:0], v3966[21:0], v5378[28:0]); // 4.0
    wire [23:0] v5379; shift_adder #(15, 22, 1, 1, 24, -9, 0) op_5379 (v3967[14:0], v3968[21:0], v5379[23:0]); // 4.0
    wire [29:0] v5380; shift_adder #(28, 17, 1, 1, 30, 13, 0) op_5380 (v3293[27:0], v3397[16:0], v5380[29:0]); // 4.0
    wire [24:0] v5381; shift_adder #(15, 24, 1, 1, 25, -9, 0) op_5381 (v3902[14:0], v3969[23:0], v5381[24:0]); // 4.0
    wire [27:0] v5382; shift_adder #(24, 26, 1, 1, 28, -3, 0) op_5382 (v3970[23:0], v3855[25:0], v5382[27:0]); // 4.0
    wire [16:0] v5383; shift_adder #(15, 16, 1, 1, 17, -1, 0) op_5383 (v3971[14:0], v3577[15:0], v5383[16:0]); // 4.0
    wire [22:0] v5384; shift_adder #(23, 19, 1, 1, 23, 2, 0) op_5384 (v3708[22:0], v3972[18:0], v5384[22:0]); // 4.0
    wire [18:0] v5385; shift_adder #(17, 15, 1, 1, 19, 3, 0) op_5385 (v3973[16:0], v3974[14:0], v5385[18:0]); // 4.0
    wire [20:0] v5386; shift_adder #(14, 21, 1, 1, 21, -4, 0) op_5386 (v3975[13:0], v3751[20:0], v5386[20:0]); // 4.0
    wire [25:0] v5387; shift_adder #(25, 13, 1, 1, 26, 11, 0) op_5387 (v3976[24:0], v3356[12:0], v5387[25:0]); // 4.0
    wire [20:0] v5388; shift_adder #(16, 20, 1, 1, 21, -5, 0) op_5388 (v3977[15:0], v3924[19:0], v5388[20:0]); // 4.0
    wire [16:0] v5389; shift_adder #(16, 15, 1, 1, 17, 1, 0) op_5389 (v3978[15:0], v2958[14:0], v5389[16:0]); // 4.0
    wire [24:0] v5390; shift_adder #(23, 24, 1, 1, 25, -1, 0) op_5390 (v2714[22:0], v3979[23:0], v5390[24:0]); // 4.0
    wire [23:0] v5391; shift_adder #(22, 15, 1, 1, 24, 9, 0) op_5391 (v3449[21:0], v3980[14:0], v5391[23:0]); // 4.0
    wire [19:0] v5392; shift_adder #(18, 15, 1, 1, 20, 4, 0) op_5392 (v3981[17:0], v2982[14:0], v5392[19:0]); // 4.0
    wire [27:0] v5393; shift_adder #(27, 17, 1, 1, 28, 11, 0) op_5393 (v3769[26:0], v2768[16:0], v5393[27:0]); // 4.0
    wire [25:0] v5394; shift_adder #(15, 26, 1, 1, 26, -10, 0) op_5394 (v3982[14:0], v3983[25:0], v5394[25:0]); // 4.0
    wire [23:0] v5395; shift_adder #(23, 19, 1, 1, 24, 5, 0) op_5395 (v3161[22:0], v3984[18:0], v5395[23:0]); // 4.0
    wire [24:0] v5396; shift_adder #(23, 25, 1, 1, 25, -1, 0) op_5396 (v3985[22:0], v3770[24:0], v5396[24:0]); // 4.0
    wire [31:0] v5397; shift_adder #(31, 27, 1, 1, 32, 5, 0) op_5397 (v3986[30:0], v3987[26:0], v5397[31:0]); // 4.0
    wire [34:0] v5398; shift_adder #(19, 35, 1, 1, 35, -14, 0) op_5398 (v3988[18:0], v3989[34:0], v5398[34:0]); // 4.0
    wire [36:0] v5399; shift_adder #(25, 36, 1, 1, 37, -10, 0) op_5399 (v3990[24:0], v3991[35:0], v5399[36:0]); // 4.0
    wire [17:0] v5400; shift_adder #(17, 15, 1, 1, 18, 1, 0) op_5400 (v3992[16:0], v3334[14:0], v5400[17:0]); // 4.0
    wire [13:0] v5401; shift_adder #(13, 13, 1, 1, 14, 0, 0) op_5401 (v3993[12:0], v2836[12:0], v5401[13:0]); // 4.0
    wire [14:0] v5402; shift_adder #(14, 14, 1, 1, 15, 1, 0) op_5402 (v3994[13:0], v3995[13:0], v5402[14:0]); // 4.0
    wire [32:0] v5403; shift_adder #(32, 32, 1, 1, 33, 0, 0) op_5403 (v3996[31:0], v3997[31:0], v5403[32:0]); // 4.0
    wire [35:0] v5404; shift_adder #(17, 35, 1, 1, 36, -19, 0) op_5404 (v3998[16:0], v3999[34:0], v5404[35:0]); // 4.0
    wire [37:0] v5405; shift_adder #(18, 37, 1, 1, 38, -19, 0) op_5405 (v4000[17:0], v4001[36:0], v5405[37:0]); // 4.0
    wire [13:0] v5406; shift_adder #(13, 12, 1, 1, 14, 0, 0) op_5406 (v4002[12:0], v3595[11:0], v5406[13:0]); // 4.0
    wire [20:0] v5407; shift_adder #(20, 19, 1, 1, 21, 1, 0) op_5407 (v3465[19:0], v4003[18:0], v5407[20:0]); // 4.0
    wire [21:0] v5408; shift_adder #(20, 22, 1, 1, 22, -1, 0) op_5408 (v2951[19:0], v4004[21:0], v5408[21:0]); // 4.0
    wire [18:0] v5409; shift_adder #(15, 17, 1, 1, 19, -3, 0) op_5409 (v4005[14:0], v4006[16:0], v5409[18:0]); // 4.0
    wire [20:0] v5410; shift_adder #(19, 21, 1, 1, 21, -1, 0) op_5410 (v4007[18:0], v3166[20:0], v5410[20:0]); // 4.0
    wire [20:0] v5411; shift_adder #(17, 20, 1, 1, 21, -3, 0) op_5411 (v3872[16:0], v2830[19:0], v5411[20:0]); // 4.0
    wire [17:0] v5412; shift_adder #(17, 16, 1, 1, 18, 1, 0) op_5412 (v4008[16:0], v4009[15:0], v5412[17:0]); // 4.0
    wire [16:0] v5413; shift_adder #(14, 15, 1, 1, 17, -2, 0) op_5413 (v4010[13:0], v4011[14:0], v5413[16:0]); // 4.0
    wire [17:0] v5414; shift_adder #(17, 17, 1, 1, 18, 1, 0) op_5414 (v3747[16:0], v4012[16:0], v5414[17:0]); // 4.0
    wire [18:0] v5415; shift_adder #(17, 14, 1, 1, 19, 4, 0) op_5415 (v4013[16:0], v2817[13:0], v5415[18:0]); // 4.0
    wire [17:0] v5416; shift_adder #(14, 16, 1, 1, 18, -3, 0) op_5416 (v3515[13:0], v4014[15:0], v5416[17:0]); // 4.0
    wire [33:0] v5417; shift_adder #(24, 32, 1, 1, 34, -9, 0) op_5417 (v4015[23:0], v2867[31:0], v5417[33:0]); // 4.0
    wire [21:0] v5418; shift_adder #(22, 21, 1, 1, 22, 0, 0) op_5418 (v3819[21:0], v3876[20:0], v5418[21:0]); // 4.0
    wire [27:0] v5419; shift_adder #(28, 20, 1, 1, 28, 7, 0) op_5419 (v3806[27:0], v4016[19:0], v5419[27:0]); // 4.0
    wire [27:0] v5420; shift_adder #(23, 27, 1, 1, 28, -4, 0) op_5420 (v3534[22:0], v2823[26:0], v5420[27:0]); // 4.0
    wire [27:0] v5421; shift_adder #(28, 15, 1, 1, 28, 12, 0) op_5421 (v2821[27:0], v4017[14:0], v5421[27:0]); // 4.0
    wire [18:0] v5422; shift_adder #(19, 17, 1, 1, 19, 0, 0) op_5422 (v4018[18:0], v4019[16:0], v5422[18:0]); // 4.0
    wire [18:0] v5423; shift_adder #(18, 15, 1, 1, 19, 3, 0) op_5423 (v4020[17:0], v4021[14:0], v5423[18:0]); // 4.0
    wire [23:0] v5424; shift_adder #(17, 24, 1, 1, 24, -4, 0) op_5424 (v3265[16:0], v3104[23:0], v5424[23:0]); // 4.0
    wire [20:0] v5425; shift_adder #(20, 18, 1, 1, 21, 1, 0) op_5425 (v4022[19:0], v4023[17:0], v5425[20:0]); // 4.0
    wire [26:0] v5426; shift_adder #(17, 24, 1, 1, 27, -10, 1) op_5426 (v615[16:0], v2527[23:0], v5426[26:0]); // 4.0
    wire [23:0] v5427; shift_adder #(20, 23, 1, 1, 24, -4, 0) op_5427 (v4024[19:0], v3210[22:0], v5427[23:0]); // 4.0
    wire [22:0] v5428; shift_adder #(14, 23, 1, 1, 23, -5, 0) op_5428 (v3459[13:0], v4025[22:0], v5428[22:0]); // 4.0
    wire [14:0] v5429; shift_adder #(14, 14, 1, 1, 15, 0, 0) op_5429 (v4026[13:0], v3853[13:0], v5429[14:0]); // 4.0
    wire [26:0] v5430; shift_adder #(25, 16, 1, 1, 27, 10, 0) op_5430 (v3670[24:0], v4027[15:0], v5430[26:0]); // 4.0
    wire [26:0] v5431; shift_adder #(14, 26, 1, 1, 27, -10, 0) op_5431 (v4028[13:0], v4029[25:0], v5431[26:0]); // 4.0
    wire [24:0] v5432; shift_adder #(24, 24, 1, 1, 25, 0, 0) op_5432 (v4030[23:0], v2781[23:0], v5432[24:0]); // 4.0
    wire [17:0] v5433; shift_adder #(16, 13, 1, 1, 18, 4, 0) op_5433 (v3920[15:0], v4031[12:0], v5433[17:0]); // 4.0
    wire [22:0] v5434; shift_adder #(16, 22, 1, 1, 23, -5, 0) op_5434 (v4032[15:0], v4033[21:0], v5434[22:0]); // 4.0
    wire [26:0] v5435; shift_adder #(27, 24, 1, 1, 27, 2, 0) op_5435 (v4034[26:0], v4035[23:0], v5435[26:0]); // 4.0
    wire [28:0] v5436; shift_adder #(28, 28, 1, 1, 29, 0, 0) op_5436 (v4036[27:0], v3325[27:0], v5436[28:0]); // 4.0
    wire [19:0] v5437; shift_adder #(19, 16, 1, 1, 20, 3, 0) op_5437 (v4003[18:0], v4037[15:0], v5437[19:0]); // 4.0
    wire [31:0] v5438; shift_adder #(19, 31, 1, 1, 32, -11, 0) op_5438 (v3470[18:0], v2889[30:0], v5438[31:0]); // 4.0
    wire [24:0] v5439; shift_adder #(25, 20, 1, 1, 25, 4, 0) op_5439 (v4038[24:0], v3785[19:0], v5439[24:0]); // 4.0
    wire [30:0] v5440; shift_adder #(30, 18, 1, 1, 31, 12, 0) op_5440 (v4039[29:0], v4040[17:0], v5440[30:0]); // 4.0
    wire [38:0] v5441; shift_adder #(37, 38, 1, 1, 39, -1, 0) op_5441 (v4041[36:0], v4042[37:0], v5441[38:0]); // 4.0
    wire [40:0] v5442; shift_adder #(25, 40, 1, 1, 41, -15, 0) op_5442 (v4043[24:0], v4044[39:0], v5442[40:0]); // 4.0
    wire [16:0] v5443; shift_adder #(16, 14, 1, 1, 17, -1, 0) op_5443 (v4045[15:0], v4046[13:0], v5443[16:0]); // 4.0
    wire [15:0] v5444; shift_adder #(15, 14, 1, 1, 16, -1, 0) op_5444 (v4047[14:0], v4048[13:0], v5444[15:0]); // 4.0
    wire [18:0] v5445; shift_adder #(18, 16, 1, 1, 19, 2, 0) op_5445 (v3483[17:0], v4049[15:0], v5445[18:0]); // 4.0
    wire [17:0] v5446; shift_adder #(14, 17, 1, 1, 18, -3, 0) op_5446 (v3768[13:0], v4050[16:0], v5446[17:0]); // 4.0
    wire [18:0] v5447; shift_adder #(17, 18, 1, 1, 19, -1, 0) op_5447 (v3794[16:0], v4051[17:0], v5447[18:0]); // 4.0
    wire [16:0] v5448; shift_adder #(16, 14, 1, 1, 17, 2, 0) op_5448 (v4052[15:0], v2871[13:0], v5448[16:0]); // 4.0
    wire [17:0] v5449; shift_adder #(16, 17, 1, 1, 18, 0, 0) op_5449 (v4053[15:0], v4054[16:0], v5449[17:0]); // 4.0
    wire [27:0] v5450; shift_adder #(18, 25, 1, 1, 28, -10, 0) op_5450 (v4055[17:0], v3672[24:0], v5450[27:0]); // 4.0
    wire [34:0] v5451; shift_adder #(31, 34, 1, 1, 35, -4, 0) op_5451 (v4056[30:0], v3492[33:0], v5451[34:0]); // 4.0
    wire [33:0] v5452; shift_adder #(34, 24, 1, 1, 34, 8, 0) op_5452 (v4057[33:0], v4058[23:0], v5452[33:0]); // 4.0
    wire [24:0] v5453; shift_adder #(24, 17, 1, 1, 25, 7, 0) op_5453 (v2519[23:0], v4059[16:0], v5453[24:0]); // 4.0
    wire [34:0] v5454; shift_adder #(34, 18, 1, 1, 35, 16, 0) op_5454 (v2874[33:0], v4023[17:0], v5454[34:0]); // 4.0
    wire [32:0] v5455; shift_adder #(15, 32, 1, 1, 33, -17, 0) op_5455 (v4060[14:0], v4061[31:0], v5455[32:0]); // 4.0
    wire [15:0] v5456; shift_adder #(16, 13, 1, 1, 16, 1, 0) op_5456 (v4062[15:0], v4063[12:0], v5456[15:0]); // 4.0
    wire [27:0] v5457; shift_adder #(10, 16, 1, 1, 28, 12, 1) op_5457 (v549[9:0], v4064[15:0], v5457[27:0]); // 4.0
    wire [29:0] v5458; shift_adder #(22, 29, 1, 1, 30, -7, 0) op_5458 (v3050[21:0], v4065[28:0], v5458[29:0]); // 4.0
    wire [25:0] v5459; shift_adder #(16, 25, 1, 1, 26, -8, 0) op_5459 (v3865[15:0], v3583[24:0], v5459[25:0]); // 4.0
    wire [30:0] v5460; shift_adder #(28, 31, 1, 1, 31, 0, 0) op_5460 (v4066[27:0], v2777[30:0], v5460[30:0]); // 4.0
    wire [27:0] v5461; shift_adder #(28, 23, 1, 1, 28, 2, 0) op_5461 (v4067[27:0], v4068[22:0], v5461[27:0]); // 4.0
    wire [18:0] v5462; shift_adder #(18, 18, 1, 1, 19, 0, 0) op_5462 (v3904[17:0], v4069[17:0], v5462[18:0]); // 4.0
    wire [21:0] v5463; shift_adder #(20, 20, 1, 1, 22, -2, 0) op_5463 (v4070[19:0], v4071[19:0], v5463[21:0]); // 4.0
    wire [15:0] v5464; shift_adder #(13, 14, 1, 1, 16, -3, 0) op_5464 (v2944[12:0], v4072[13:0], v5464[15:0]); // 4.0
    wire [20:0] v5465; shift_adder #(20, 15, 1, 1, 21, 5, 0) op_5465 (v3532[19:0], v4073[14:0], v5465[20:0]); // 4.0
    wire [15:0] v5466; shift_adder #(13, 14, 1, 1, 16, 1, 0) op_5466 (v4074[12:0], v4075[13:0], v5466[15:0]); // 4.0
    wire [18:0] v5467; shift_adder #(17, 14, 1, 1, 19, 4, 0) op_5467 (v4076[16:0], v4077[13:0], v5467[18:0]); // 4.0
    wire [20:0] v5468; shift_adder #(15, 21, 1, 1, 21, -3, 0) op_5468 (v4078[14:0], v4079[20:0], v5468[20:0]); // 4.0
    wire [16:0] v5469; shift_adder #(15, 16, 1, 1, 17, 0, 0) op_5469 (v4080[14:0], v2513[15:0], v5469[16:0]); // 4.0
    wire [20:0] v5470; shift_adder #(18, 19, 1, 1, 21, -2, 0) op_5470 (v4081[17:0], v4082[18:0], v5470[20:0]); // 4.0
    wire [24:0] v5471; shift_adder #(22, 18, 1, 1, 25, 7, 0) op_5471 (v3037[21:0], v4083[17:0], v5471[24:0]); // 4.0
    wire [20:0] v5472; shift_adder #(20, 15, 1, 1, 21, 5, 0) op_5472 (v4022[19:0], v3443[14:0], v5472[20:0]); // 4.0
    wire [32:0] v5473; shift_adder #(32, 18, 1, 1, 33, 14, 0) op_5473 (v4084[31:0], v3631[17:0], v5473[32:0]); // 4.0
    wire [25:0] v5474; shift_adder #(14, 25, 1, 1, 26, -12, 0) op_5474 (v4085[13:0], v3680[24:0], v5474[25:0]); // 4.0
    wire [15:0] v5475; shift_adder #(14, 14, 1, 1, 16, -1, 0) op_5475 (v4086[13:0], v4087[13:0], v5475[15:0]); // 4.0
    wire [25:0] v5476; shift_adder #(25, 21, 1, 1, 26, 4, 0) op_5476 (v4088[24:0], v3873[20:0], v5476[25:0]); // 4.0
    wire [29:0] v5477; shift_adder #(29, 13, 1, 1, 30, 16, 0) op_5477 (v4089[28:0], v3151[12:0], v5477[29:0]); // 4.0
    wire [23:0] v5478; shift_adder #(17, 23, 1, 1, 24, -6, 0) op_5478 (v4090[16:0], v4091[22:0], v5478[23:0]); // 4.0
    wire [33:0] v5479; shift_adder #(26, 33, 1, 1, 34, -7, 0) op_5479 (v4092[25:0], v4093[32:0], v5479[33:0]); // 4.0
    wire [27:0] v5480; shift_adder #(27, 20, 1, 1, 28, 6, 0) op_5480 (v4094[26:0], v3802[19:0], v5480[27:0]); // 4.0
    wire [36:0] v5481; shift_adder #(35, 19, 1, 1, 37, 17, 0) op_5481 (v4095[34:0], v3753[18:0], v5481[36:0]); // 4.0
    wire [37:0] v5482; shift_adder #(16, 14, 1, 1, 38, 24, 1) op_5482 (v4096[15:0], v2304[13:0], v5482[37:0]); // 4.0
    wire [36:0] v5483; shift_adder #(37, 14, 1, 1, 37, 1, 1) op_5483 (v4097[36:0], v4098[13:0], v5483[36:0]); // 4.0
    wire [17:0] v5484; shift_adder #(17, 15, 1, 1, 18, 1, 0) op_5484 (v4099[16:0], v4100[14:0], v5484[17:0]); // 4.0
    wire [16:0] v5485; shift_adder #(16, 14, 1, 1, 17, 2, 0) op_5485 (v4101[15:0], v2719[13:0], v5485[16:0]); // 4.0
    wire [36:0] v5486; shift_adder #(13, 36, 1, 1, 37, -22, 0) op_5486 (v4102[12:0], v4103[35:0], v5486[36:0]); // 4.0
    wire [18:0] v5487; shift_adder #(19, 14, 1, 1, 19, 2, 0) op_5487 (v3988[18:0], v2552[13:0], v5487[18:0]); // 4.0
    wire [19:0] v5488; shift_adder #(19, 12, 1, 1, 20, 5, 0) op_5488 (v4104[18:0], v3174[11:0], v5488[19:0]); // 4.0
    wire [17:0] v5489; shift_adder #(15, 17, 1, 1, 18, -1, 0) op_5489 (v3032[14:0], v4105[16:0], v5489[17:0]); // 4.0
    wire [16:0] v5490; shift_adder #(16, 14, 1, 1, 17, 2, 0) op_5490 (v4106[15:0], v3711[13:0], v5490[16:0]); // 4.0
    wire [16:0] v5491; shift_adder #(16, 16, 1, 1, 17, 0, 0) op_5491 (v3091[15:0], v2918[15:0], v5491[16:0]); // 4.0
    wire [30:0] v5492; shift_adder #(30, 16, 1, 1, 31, 13, 0) op_5492 (v4107[29:0], v4108[15:0], v5492[30:0]); // 4.0
    wire [26:0] v5493; shift_adder #(26, 25, 1, 1, 27, 0, 0) op_5493 (v4109[25:0], v4110[24:0], v5493[26:0]); // 4.0
    wire [26:0] v5494; shift_adder #(25, 22, 1, 1, 27, 4, 0) op_5494 (v4111[24:0], v3808[21:0], v5494[26:0]); // 4.0
    wire [18:0] v5495; shift_adder #(19, 14, 1, 1, 19, 3, 0) op_5495 (v3221[18:0], v4112[13:0], v5495[18:0]); // 4.0
    wire [26:0] v5496; shift_adder #(20, 25, 1, 1, 27, -7, 0) op_5496 (v3178[19:0], v4113[24:0], v5496[26:0]); // 4.0
    wire [26:0] v5497; shift_adder #(22, 26, 1, 1, 27, -5, 0) op_5497 (v4114[21:0], v4115[25:0], v5497[26:0]); // 4.0
    wire [15:0] v5498; shift_adder #(14, 15, 1, 1, 16, -2, 0) op_5498 (v4116[13:0], v4117[14:0], v5498[15:0]); // 4.0
    wire [23:0] v5499; shift_adder #(24, 22, 1, 1, 24, 1, 0) op_5499 (v4118[23:0], v4119[21:0], v5499[23:0]); // 4.0
    wire [21:0] v5500; shift_adder #(22, 20, 1, 1, 22, 0, 0) op_5500 (v4120[21:0], v4121[19:0], v5500[21:0]); // 4.0
    wire [20:0] v5501; shift_adder #(20, 15, 1, 1, 21, 6, 0) op_5501 (v4122[19:0], v4123[14:0], v5501[20:0]); // 4.0
    wire [20:0] v5502; shift_adder #(18, 20, 1, 1, 21, -2, 0) op_5502 (v4124[17:0], v4125[19:0], v5502[20:0]); // 4.0
    wire [18:0] v5503; shift_adder #(13, 18, 1, 1, 19, -4, 0) op_5503 (v4126[12:0], v4127[17:0], v5503[18:0]); // 4.0
    wire [17:0] v5504; shift_adder #(16, 17, 1, 1, 18, 0, 0) op_5504 (v4128[15:0], v4129[16:0], v5504[17:0]); // 4.0
    wire [16:0] v5505; shift_adder #(16, 15, 1, 1, 17, 1, 0) op_5505 (v3915[15:0], v4130[14:0], v5505[16:0]); // 4.0
    wire [21:0] v5506; shift_adder #(20, 22, 1, 1, 22, -1, 0) op_5506 (v4131[19:0], v3501[21:0], v5506[21:0]); // 4.0
    wire [18:0] v5507; shift_adder #(18, 18, 1, 1, 19, 0, 0) op_5507 (v4132[17:0], v3074[17:0], v5507[18:0]); // 4.0
    wire [17:0] v5508; shift_adder #(13, 17, 1, 1, 18, -3, 0) op_5508 (v3093[12:0], v4133[16:0], v5508[17:0]); // 4.0
    wire [21:0] v5509; shift_adder #(18, 22, 1, 1, 22, -1, 0) op_5509 (v4040[17:0], v3224[21:0], v5509[21:0]); // 4.0
    wire [23:0] v5510; shift_adder #(23, 19, 1, 1, 24, 5, 0) op_5510 (v4134[22:0], v4135[18:0], v5510[23:0]); // 4.0
    wire [23:0] v5511; shift_adder #(23, 24, 1, 1, 24, 0, 0) op_5511 (v4136[22:0], v3121[23:0], v5511[23:0]); // 4.0
    wire [24:0] v5512; shift_adder #(24, 17, 1, 1, 25, 7, 0) op_5512 (v3653[23:0], v4137[16:0], v5512[24:0]); // 4.0
    wire [31:0] v5513; shift_adder #(9, 32, 1, 1, 32, -21, 0) op_5513 (v490[8:0], v4138[31:0], v5513[31:0]); // 4.0
    wire [20:0] v5514; shift_adder #(14, 20, 1, 1, 21, -4, 0) op_5514 (v3136[13:0], v4139[19:0], v5514[20:0]); // 4.0
    wire [33:0] v5515; shift_adder #(33, 14, 1, 1, 34, 20, 0) op_5515 (v4140[32:0], v4141[13:0], v5515[33:0]); // 4.0
    wire [38:0] v5516; shift_adder #(24, 38, 1, 1, 39, -13, 0) op_5516 (v4142[23:0], v4143[37:0], v5516[38:0]); // 4.0
    wire [16:0] v5517; shift_adder #(14, 14, 1, 1, 17, -2, 0) op_5517 (v2586[13:0], v4144[13:0], v5517[16:0]); // 4.0
    wire [20:0] v5518; shift_adder #(21, 20, 1, 1, 21, 0, 0) op_5518 (v3051[20:0], v3798[19:0], v5518[20:0]); // 4.0
    wire [22:0] v5519; shift_adder #(13, 22, 1, 1, 23, -10, 0) op_5519 (v4145[12:0], v2604[21:0], v5519[22:0]); // 4.0
    wire [19:0] v5520; shift_adder #(15, 19, 1, 1, 20, -3, 0) op_5520 (v4146[14:0], v4147[18:0], v5520[19:0]); // 4.0
    wire [18:0] v5521; shift_adder #(19, 15, 1, 1, 19, 3, 0) op_5521 (v4148[18:0], v2765[14:0], v5521[18:0]); // 4.0
    wire [31:0] v5522; shift_adder #(31, 20, 1, 1, 32, 12, 0) op_5522 (v2741[30:0], v2723[19:0], v5522[31:0]); // 4.0
    wire [15:0] v5523; shift_adder #(14, 13, 1, 1, 16, 2, 0) op_5523 (v4149[13:0], v4150[12:0], v5523[15:0]); // 4.0
    wire [15:0] v5524; shift_adder #(14, 15, 1, 1, 16, -1, 0) op_5524 (v4151[13:0], v2622[14:0], v5524[15:0]); // 4.0
    wire [20:0] v5525; shift_adder #(13, 20, 1, 1, 21, -7, 0) op_5525 (v3888[12:0], v4153[19:0], v5525[20:0]); // 4.0
    wire [39:0] v5526; shift_adder #(40, 16, 1, 1, 40, 23, 0) op_5526 (v4154[39:0], v3207[15:0], v5526[39:0]); // 4.0
    wire [35:0] v5527; shift_adder #(18, 14, 1, 1, 36, -18, 1) op_5527 (v4051[17:0], v4155[13:0], v5527[35:0]); // 4.0
    wire [23:0] v5528; shift_adder #(15, 24, 1, 1, 24, -8, 0) op_5528 (v2996[14:0], v3821[23:0], v5528[23:0]); // 4.0
    wire [31:0] v5529; shift_adder #(17, 30, 1, 1, 32, -14, 0) op_5529 (v4156[16:0], v4157[29:0], v5529[31:0]); // 4.0
    wire [27:0] v5530; shift_adder #(20, 27, 1, 1, 28, -7, 0) op_5530 (v4158[19:0], v4159[26:0], v5530[27:0]); // 4.0
    wire [26:0] v5531; shift_adder #(26, 20, 1, 1, 27, 6, 0) op_5531 (v4160[25:0], v2873[19:0], v5531[26:0]); // 4.0
    wire [32:0] v5532; shift_adder #(15, 32, 1, 1, 33, -17, 0) op_5532 (v3939[14:0], v3996[31:0], v5532[32:0]); // 4.0
    wire [30:0] v5533; shift_adder #(24, 31, 1, 1, 31, -5, 0) op_5533 (v3079[23:0], v4161[30:0], v5533[30:0]); // 4.0
    wire [15:0] v5534; shift_adder #(15, 15, 1, 1, 16, 1, 0) op_5534 (v4162[14:0], v4163[14:0], v5534[15:0]); // 4.0
    wire [24:0] v5535; shift_adder #(25, 14, 1, 1, 25, 8, 0) op_5535 (v4164[24:0], v4048[13:0], v5535[24:0]); // 4.0
    wire [28:0] v5536; shift_adder #(26, 28, 1, 1, 29, -2, 0) op_5536 (v4165[25:0], v2789[27:0], v5536[28:0]); // 4.0
    wire [18:0] v5537; shift_adder #(18, 14, 1, 1, 19, 3, 0) op_5537 (v4166[17:0], v2991[13:0], v5537[18:0]); // 4.0
    wire [23:0] v5538; shift_adder #(24, 17, 1, 1, 24, 4, 0) op_5538 (v3060[23:0], v4167[16:0], v5538[23:0]); // 4.0
    wire [25:0] v5539; shift_adder #(26, 22, 1, 1, 26, 2, 0) op_5539 (v4168[25:0], v4169[21:0], v5539[25:0]); // 4.0
    wire [17:0] v5540; shift_adder #(18, 16, 1, 1, 18, 1, 0) op_5540 (v4170[17:0], v4171[15:0], v5540[17:0]); // 4.0
    wire [22:0] v5541; shift_adder #(21, 14, 1, 1, 23, 9, 0) op_5541 (v4172[20:0], v4173[13:0], v5541[22:0]); // 4.0
    wire [23:0] v5542; shift_adder #(14, 24, 1, 1, 24, -8, 0) op_5542 (v4174[13:0], v4175[23:0], v5542[23:0]); // 4.0
    wire [22:0] v5543; shift_adder #(22, 14, 1, 1, 23, 9, 0) op_5543 (v4176[21:0], v4177[13:0], v5543[22:0]); // 4.0
    wire [28:0] v5544; shift_adder #(28, 22, 1, 1, 29, 6, 0) op_5544 (v4178[27:0], v4179[21:0], v5544[28:0]); // 4.0
    wire [28:0] v5545; shift_adder #(19, 26, 1, 1, 29, -10, 0) op_5545 (v3879[18:0], v4165[25:0], v5545[28:0]); // 4.0
    wire [17:0] v5546; shift_adder #(15, 16, 1, 1, 18, -2, 0) op_5546 (v2710[14:0], v2566[15:0], v5546[17:0]); // 4.0
    wire [18:0] v5547; shift_adder #(16, 17, 1, 1, 19, -3, 0) op_5547 (v4180[15:0], v3231[16:0], v5547[18:0]); // 4.0
    wire [26:0] v5548; shift_adder #(26, 19, 1, 1, 27, 8, 0) op_5548 (v2632[25:0], v4181[18:0], v5548[26:0]); // 4.0
    wire [26:0] v5549; shift_adder #(16, 25, 1, 1, 27, -11, 0) op_5549 (v3437[15:0], v3414[24:0], v5549[26:0]); // 4.0
    wire [24:0] v5550; shift_adder #(14, 24, 1, 1, 25, -10, 0) op_5550 (v3028[13:0], v3052[23:0], v5550[24:0]); // 4.0
    wire [24:0] v5551; shift_adder #(24, 12, 1, 1, 25, 11, 0) op_5551 (v4182[23:0], v2733[11:0], v5551[24:0]); // 4.0
    wire [28:0] v5552; shift_adder #(28, 14, 1, 1, 29, 14, 0) op_5552 (v4183[27:0], v4184[13:0], v5552[28:0]); // 4.0
    wire [26:0] v5553; shift_adder #(27, 17, 1, 1, 27, 8, 0) op_5553 (v4185[26:0], v4186[16:0], v5553[26:0]); // 4.0
    wire [29:0] v5554; shift_adder #(29, 14, 1, 1, 30, 15, 0) op_5554 (v4089[28:0], v4187[13:0], v5554[29:0]); // 4.0
    wire [22:0] v5555; shift_adder #(22, 16, 1, 1, 23, 6, 0) op_5555 (v3757[21:0], v3765[15:0], v5555[22:0]); // 4.0
    wire [26:0] v5556; shift_adder #(15, 26, 1, 1, 27, -11, 0) op_5556 (v4188[14:0], v3703[25:0], v5556[26:0]); // 4.0
    wire [19:0] v5557; shift_adder #(17, 20, 1, 1, 20, -1, 0) op_5557 (v4189[16:0], v3487[19:0], v5557[19:0]); // 4.0
    wire [32:0] v5558; shift_adder #(32, 18, 1, 1, 33, 15, 0) op_5558 (v4190[31:0], v4191[17:0], v5558[32:0]); // 4.0
    wire [35:0] v5559; shift_adder #(16, 35, 1, 1, 36, -18, 0) op_5559 (v4192[15:0], v4193[34:0], v5559[35:0]); // 4.0
    wire [19:0] v5560; shift_adder #(19, 15, 1, 1, 20, 4, 0) op_5560 (v4194[18:0], v4195[14:0], v5560[19:0]); // 4.0
    wire [20:0] v5561; shift_adder #(18, 19, 1, 1, 21, 2, 0) op_5561 (v3523[17:0], v4196[18:0], v5561[20:0]); // 4.0
    wire [34:0] v5562; shift_adder #(16, 33, 1, 1, 35, -18, 0) op_5562 (v4197[15:0], v4198[32:0], v5562[34:0]); // 4.0
    wire [28:0] v5563; shift_adder #(19, 27, 1, 1, 29, -10, 0) op_5563 (v2999[18:0], v3959[26:0], v5563[28:0]); // 4.0
    wire [39:0] v5564; shift_adder #(16, 40, 1, 1, 40, -22, 0) op_5564 (v2970[15:0], v4199[39:0], v5564[39:0]); // 4.0
    wire [17:0] v5565; shift_adder #(17, 14, 1, 1, 18, 4, 0) op_5565 (v4200[16:0], v4201[13:0], v5565[17:0]); // 4.0
    wire [38:0] v5566; shift_adder #(34, 38, 1, 1, 39, -4, 0) op_5566 (v4202[33:0], v4203[37:0], v5566[38:0]); // 4.0
    wire [14:0] v5567; shift_adder #(14, 15, 1, 1, 15, 0, 0) op_5567 (v4204[13:0], v4205[14:0], v5567[14:0]); // 4.0
    wire [14:0] v5568; shift_adder #(13, 12, 1, 1, 15, -1, 0) op_5568 (v3993[12:0], v4206[11:0], v5568[14:0]); // 4.0
    wire [21:0] v5569; shift_adder #(21, 16, 1, 1, 22, 3, 0) op_5569 (v3522[20:0], v4207[15:0], v5569[21:0]); // 4.0
    wire [25:0] v5570; shift_adder #(25, 19, 1, 1, 26, 4, 0) op_5570 (v4208[24:0], v4209[18:0], v5570[25:0]); // 4.0
    wire [22:0] v5571; shift_adder #(14, 21, 1, 1, 23, -8, 0) op_5571 (v4210[13:0], v4211[20:0], v5571[22:0]); // 4.0
    wire [19:0] v5572; shift_adder #(18, 19, 1, 1, 20, -1, 0) op_5572 (v4212[17:0], v4213[18:0], v5572[19:0]); // 4.0
    wire [19:0] v5573; shift_adder #(18, 19, 1, 1, 20, -2, 0) op_5573 (v4214[17:0], v4215[18:0], v5573[19:0]); // 4.0
    wire [15:0] v5574; shift_adder #(13, 15, 1, 1, 16, -1, 0) op_5574 (v4216[12:0], v4217[14:0], v5574[15:0]); // 4.0
    wire [15:0] v5575; shift_adder #(14, 14, 1, 1, 16, -1, 0) op_5575 (v4218[13:0], v4219[13:0], v5575[15:0]); // 4.0
    wire [16:0] v5576; shift_adder #(16, 16, 1, 1, 17, 0, 0) op_5576 (v3205[15:0], v4220[15:0], v5576[16:0]); // 4.0
    wire [19:0] v5577; shift_adder #(18, 19, 1, 1, 20, 1, 0) op_5577 (v4221[17:0], v4222[18:0], v5577[19:0]); // 4.0
    wire [21:0] v5578; shift_adder #(13, 22, 1, 1, 22, -7, 0) op_5578 (v4223[12:0], v4120[21:0], v5578[21:0]); // 4.0
    wire [20:0] v5579; shift_adder #(16, 21, 1, 1, 21, -4, 0) op_5579 (v4224[15:0], v4225[20:0], v5579[20:0]); // 4.0
    wire [21:0] v5580; shift_adder #(14, 21, 1, 1, 22, -7, 0) op_5580 (v2664[13:0], v4226[20:0], v5580[21:0]); // 4.0
    wire [22:0] v5581; shift_adder #(22, 20, 1, 1, 23, 3, 0) op_5581 (v4179[21:0], v3962[19:0], v5581[22:0]); // 4.0
    wire [23:0] v5582; shift_adder #(23, 18, 1, 1, 24, 5, 0) op_5582 (v4227[22:0], v4228[17:0], v5582[23:0]); // 4.0
    wire [20:0] v5583; shift_adder #(19, 20, 1, 1, 21, 0, 0) op_5583 (v4229[18:0], v4230[19:0], v5583[20:0]); // 4.0
    wire [27:0] v5584; shift_adder #(26, 21, 1, 1, 28, 6, 0) op_5584 (v3866[25:0], v2846[20:0], v5584[27:0]); // 4.0
    wire [28:0] v5585; shift_adder #(18, 28, 1, 1, 29, -11, 0) op_5585 (v4231[17:0], v3563[27:0], v5585[28:0]); // 4.0
    wire [18:0] v5586; shift_adder #(15, 18, 1, 1, 19, -1, 0) op_5586 (v4232[14:0], v4233[17:0], v5586[18:0]); // 4.0
    wire [26:0] v5587; shift_adder #(14, 27, 1, 1, 27, -12, 0) op_5587 (v4234[13:0], v2736[26:0], v5587[26:0]); // 4.0
    wire [27:0] v5588; shift_adder #(26, 28, 1, 1, 28, 0, 0) op_5588 (v4235[25:0], v4236[27:0], v5588[27:0]); // 4.0
    wire [30:0] v5589; shift_adder #(8, 23, 1, 1, 31, -22, 0) op_5589 (v93[7:0], v4237[22:0], v5589[30:0]); // 4.0
    wire [15:0] v5590; shift_adder #(16, 14, 1, 1, 16, 1, 0) op_5590 (v4238[15:0], v3369[13:0], v5590[15:0]); // 4.0
    wire [20:0] v5591; shift_adder #(19, 20, 1, 1, 21, -1, 0) op_5591 (v4240[18:0], v3640[19:0], v5591[20:0]); // 4.0
    wire [18:0] v5592; shift_adder #(18, 15, 1, 1, 19, 2, 0) op_5592 (v4233[17:0], v4241[14:0], v5592[18:0]); // 4.0
    wire [24:0] v5593; shift_adder #(16, 24, 1, 1, 25, -7, 0) op_5593 (v4242[15:0], v4243[23:0], v5593[24:0]); // 4.0
    wire [35:0] v5594; shift_adder #(14, 12, 1, 1, 36, 24, 1) op_5594 (v3557[13:0], v2393[11:0], v5594[35:0]); // 4.0
    wire [37:0] v5595; shift_adder #(38, 24, 1, 1, 38, 13, 0) op_5595 (v4244[37:0], v3979[23:0], v5595[37:0]); // 4.0
    wire [28:0] v5596; shift_adder #(24, 28, 1, 1, 29, -4, 0) op_5596 (v3341[23:0], v4245[27:0], v5596[28:0]); // 4.0
    wire [15:0] v5597; shift_adder #(13, 16, 1, 1, 16, -2, 0) op_5597 (v4246[12:0], v4247[15:0], v5597[15:0]); // 4.0
    wire [14:0] v5598; shift_adder #(13, 14, 1, 1, 15, -1, 0) op_5598 (v2575[12:0], v3527[13:0], v5598[14:0]); // 4.0
    wire [15:0] v5599; shift_adder #(15, 15, 1, 1, 16, 1, 0) op_5599 (v4248[14:0], v2593[14:0], v5599[15:0]); // 4.0
    wire [15:0] v5600; shift_adder #(15, 13, 1, 1, 16, 1, 0) op_5600 (v4249[14:0], v4063[12:0], v5600[15:0]); // 4.0
    wire [33:0] v5601; shift_adder #(19, 33, 1, 1, 34, -15, 0) op_5601 (v4250[18:0], v4251[32:0], v5601[33:0]); // 4.0
    wire [31:0] v5602; shift_adder #(31, 22, 1, 1, 32, 9, 0) op_5602 (v2576[30:0], v4252[21:0], v5602[31:0]); // 4.0
    wire [21:0] v5603; shift_adder #(22, 16, 1, 1, 22, 4, 0) op_5603 (v4253[21:0], v4254[15:0], v5603[21:0]); // 4.0
    wire [27:0] v5604; shift_adder #(28, 20, 1, 1, 28, 6, 0) op_5604 (v3481[27:0], v3021[19:0], v5604[27:0]); // 4.0
    wire [25:0] v5605; shift_adder #(23, 25, 1, 1, 26, -3, 0) op_5605 (v3761[22:0], v4255[24:0], v5605[25:0]); // 4.0
    wire [26:0] v5606; shift_adder #(26, 26, 1, 1, 27, -1, 0) op_5606 (v4256[25:0], v4257[25:0], v5606[26:0]); // 4.0
    wire [25:0] v5607; shift_adder #(19, 24, 1, 1, 26, -6, 0) op_5607 (v4258[18:0], v4259[23:0], v5607[25:0]); // 4.0
    wire [22:0] v5608; shift_adder #(16, 21, 1, 1, 23, -6, 0) op_5608 (v3169[15:0], v3789[20:0], v5608[22:0]); // 4.0
    wire [16:0] v5609; shift_adder #(14, 16, 1, 1, 17, -1, 0) op_5609 (v4260[13:0], v4261[15:0], v5609[16:0]); // 4.0
    wire [25:0] v5610; shift_adder #(24, 25, 1, 1, 26, -2, 0) op_5610 (v2931[23:0], v3990[24:0], v5610[25:0]); // 4.0
    wire [20:0] v5611; shift_adder #(15, 21, 1, 1, 21, -4, 0) op_5611 (v4262[14:0], v4263[20:0], v5611[20:0]); // 4.0
    wire [22:0] v5612; shift_adder #(22, 18, 1, 1, 23, 3, 0) op_5612 (v4264[21:0], v2690[17:0], v5612[22:0]); // 4.0
    wire [23:0] v5613; shift_adder #(18, 23, 1, 1, 24, -5, 0) op_5613 (v3671[17:0], v4265[22:0], v5613[23:0]); // 4.0
    wire [19:0] v5614; shift_adder #(17, 19, 1, 1, 20, -1, 0) op_5614 (v4266[16:0], v3949[18:0], v5614[19:0]); // 4.0
    wire [19:0] v5615; shift_adder #(16, 20, 1, 1, 20, -3, 0) op_5615 (v4267[15:0], v3262[19:0], v5615[19:0]); // 4.0
    wire [21:0] v5616; shift_adder #(21, 18, 1, 1, 22, 3, 0) op_5616 (v4268[20:0], v4269[17:0], v5616[21:0]); // 4.0
    wire [25:0] v5617; shift_adder #(18, 25, 1, 1, 26, -5, 0) op_5617 (v4020[17:0], v4270[24:0], v5617[25:0]); // 4.0
    wire [29:0] v5618; shift_adder #(27, 30, 1, 1, 30, 0, 0) op_5618 (v2623[26:0], v4271[29:0], v5618[29:0]); // 4.0
    wire [29:0] v5619; shift_adder #(28, 24, 1, 1, 30, 6, 0) op_5619 (v4272[27:0], v4273[23:0], v5619[29:0]); // 4.0
    wire [28:0] v5620; shift_adder #(15, 28, 1, 1, 29, -13, 0) op_5620 (v3857[14:0], v4274[27:0], v5620[28:0]); // 4.0
    wire [22:0] v5621; shift_adder #(22, 15, 1, 1, 23, 8, 0) op_5621 (v3261[21:0], v4275[14:0], v5621[22:0]); // 4.0
    wire [22:0] v5622; shift_adder #(22, 21, 1, 1, 23, 0, 0) op_5622 (v3966[21:0], v4276[20:0], v5622[22:0]); // 4.0
    wire [19:0] v5623; shift_adder #(17, 20, 1, 1, 20, -1, 0) op_5623 (v4277[16:0], v4278[19:0], v5623[19:0]); // 4.0
    wire [25:0] v5624; shift_adder #(13, 26, 1, 1, 26, -10, 0) op_5624 (v3542[12:0], v3120[25:0], v5624[25:0]); // 4.0
    wire [23:0] v5625; shift_adder #(16, 24, 1, 1, 24, -6, 0) op_5625 (v4279[15:0], v4280[23:0], v5625[23:0]); // 4.0
    wire [18:0] v5626; shift_adder #(18, 17, 1, 1, 19, 1, 0) op_5626 (v4228[17:0], v2922[16:0], v5626[18:0]); // 4.0
    wire [22:0] v5627; shift_adder #(22, 17, 1, 1, 23, 5, 0) op_5627 (v4281[21:0], v4282[16:0], v5627[22:0]); // 4.0
    wire [17:0] v5628; shift_adder #(14, 17, 1, 1, 18, -3, 0) op_5628 (v4283[13:0], v4284[16:0], v5628[17:0]); // 4.0
    wire [14:0] v5629; shift_adder #(12, 15, 1, 1, 15, -2, 0) op_5629 (v2973[11:0], v4285[14:0], v5629[14:0]); // 4.0
    wire [38:0] v5630; shift_adder #(17, 38, 1, 1, 39, -21, 0) op_5630 (v4287[16:0], v4288[37:0], v5630[38:0]); // 4.0
    wire [20:0] v5631; shift_adder #(14, 19, 1, 1, 21, -6, 0) op_5631 (v4289[13:0], v4290[18:0], v5631[20:0]); // 4.0
    wire [18:0] v5632; shift_adder #(19, 15, 1, 1, 19, 3, 0) op_5632 (v3243[18:0], v4291[14:0], v5632[18:0]); // 4.0
    wire [20:0] v5633; shift_adder #(20, 17, 1, 1, 21, 3, 0) op_5633 (v3755[19:0], v4292[16:0], v5633[20:0]); // 4.0
    wire [17:0] v5634; shift_adder #(17, 17, 1, 1, 18, 0, 0) op_5634 (v4293[16:0], v4294[16:0], v5634[17:0]); // 4.0
    wire [41:0] v5635; shift_adder #(42, 14, 1, 1, 42, 3, 1) op_5635 (v4295[41:0], v4296[13:0], v5635[41:0]); // 4.0
    wire [18:0] v5636; shift_adder #(19, 16, 1, 1, 19, 0, 0) op_5636 (v4297[18:0], v4298[15:0], v5636[18:0]); // 4.0
    wire [15:0] v5637; shift_adder #(15, 13, 1, 1, 16, 2, 0) op_5637 (v4299[14:0], v4300[12:0], v5637[15:0]); // 4.0
    wire [16:0] v5638; shift_adder #(15, 16, 1, 1, 17, 0, 0) op_5638 (v4301[14:0], v4302[15:0], v5638[16:0]); // 4.0
    wire [22:0] v5639; shift_adder #(22, 12, 1, 1, 23, 10, 0) op_5639 (v3607[21:0], v4303[11:0], v5639[22:0]); // 4.0
    wire [32:0] v5640; shift_adder #(32, 30, 1, 1, 33, 2, 0) op_5640 (v2800[31:0], v4304[29:0], v5640[32:0]); // 4.0
    wire [18:0] v5641; shift_adder #(16, 17, 1, 1, 19, -2, 0) op_5641 (v4305[15:0], v3432[16:0], v5641[18:0]); // 4.0
    wire [23:0] v5642; shift_adder #(18, 23, 1, 1, 24, -6, 0) op_5642 (v4306[17:0], v3815[22:0], v5642[23:0]); // 4.0
    wire [29:0] v5643; shift_adder #(17, 28, 1, 1, 30, -12, 0) op_5643 (v3601[16:0], v4307[27:0], v5643[29:0]); // 4.0
    wire [28:0] v5644; shift_adder #(26, 28, 1, 1, 29, -2, 0) op_5644 (v2679[25:0], v4308[27:0], v5644[28:0]); // 4.0
    wire [22:0] v5645; shift_adder #(23, 17, 1, 1, 23, 5, 0) op_5645 (v3336[22:0], v4309[16:0], v5645[22:0]); // 4.0
    wire [29:0] v5646; shift_adder #(19, 29, 1, 1, 30, -11, 0) op_5646 (v4310[18:0], v4311[28:0], v5646[29:0]); // 4.0
    wire [27:0] v5647; shift_adder #(27, 23, 1, 1, 28, 4, 0) op_5647 (v4312[26:0], v3908[22:0], v5647[27:0]); // 4.0
    wire [24:0] v5648; shift_adder #(24, 20, 1, 1, 25, 3, 0) op_5648 (v4313[23:0], v4314[19:0], v5648[24:0]); // 4.0
    wire [26:0] v5649; shift_adder #(13, 26, 1, 1, 27, -12, 0) op_5649 (v4315[12:0], v3511[25:0], v5649[26:0]); // 4.0
    wire [17:0] v5650; shift_adder #(8, 18, 1, 1, 18, -2, 1) op_5650 (v89[7:0], v4316[17:0], v5650[17:0]); // 4.0
    wire [18:0] v5651; shift_adder #(15, 19, 1, 1, 19, -3, 0) op_5651 (v3967[14:0], v3271[18:0], v5651[18:0]); // 4.0
    wire [16:0] v5652; shift_adder #(14, 13, 1, 1, 17, 3, 0) op_5652 (v4317[13:0], v4315[12:0], v5652[16:0]); // 4.0
    wire [17:0] v5653; shift_adder #(17, 14, 1, 1, 18, 2, 0) op_5653 (v4318[16:0], v2901[13:0], v5653[17:0]); // 4.0
    wire [17:0] v5654; shift_adder #(14, 17, 1, 1, 18, -3, 0) op_5654 (v4319[13:0], v2641[16:0], v5654[17:0]); // 4.0
    wire [15:0] v5655; shift_adder #(15, 13, 1, 1, 16, 2, 0) op_5655 (v4320[14:0], v3524[12:0], v5655[15:0]); // 4.0
    wire [19:0] v5656; shift_adder #(19, 13, 1, 1, 20, 7, 0) op_5656 (v4321[18:0], v2545[12:0], v5656[19:0]); // 4.0
    wire [15:0] v5657; shift_adder #(15, 15, 1, 1, 16, 1, 0) op_5657 (v4322[14:0], v4323[14:0], v5657[15:0]); // 4.0
    wire [21:0] v5658; shift_adder #(20, 15, 1, 1, 22, 6, 0) op_5658 (v3021[19:0], v4324[14:0], v5658[21:0]); // 4.0
    wire [24:0] v5659; shift_adder #(17, 23, 1, 1, 25, -7, 0) op_5659 (v4156[16:0], v4325[22:0], v5659[24:0]); // 4.0
    wire [30:0] v5660; shift_adder #(14, 28, 1, 1, 31, -17, 0) op_5660 (v4326[13:0], v3215[27:0], v5660[30:0]); // 4.0
    wire [22:0] v5661; shift_adder #(21, 21, 1, 1, 23, -1, 0) op_5661 (v4327[20:0], v4328[20:0], v5661[22:0]); // 4.0
    wire [30:0] v5662; shift_adder #(13, 29, 1, 1, 31, -18, 0) op_5662 (v3083[12:0], v4329[28:0], v5662[30:0]); // 4.0
    wire [29:0] v5663; shift_adder #(23, 30, 1, 1, 30, -4, 0) op_5663 (v4330[22:0], v3870[29:0], v5663[29:0]); // 4.0
    wire [15:0] v5664; shift_adder #(15, 16, 1, 1, 16, 0, 0) op_5664 (v3738[14:0], v4331[15:0], v5664[15:0]); // 4.0
    wire [27:0] v5665; shift_adder #(14, 27, 1, 1, 28, -13, 0) op_5665 (v4116[13:0], v4332[26:0], v5665[27:0]); // 4.0
    wire [30:0] v5666; shift_adder #(29, 26, 1, 1, 31, 5, 0) op_5666 (v4311[28:0], v3073[25:0], v5666[30:0]); // 4.0
    wire [31:0] v5667; shift_adder #(32, 25, 1, 1, 32, 6, 0) op_5667 (v3567[31:0], v4333[24:0], v5667[31:0]); // 4.0
    wire [23:0] v5668; shift_adder #(24, 22, 1, 1, 24, 1, 0) op_5668 (v2815[23:0], v2924[21:0], v5668[23:0]); // 4.0
    wire [19:0] v5669; shift_adder #(19, 16, 1, 1, 20, 3, 0) op_5669 (v4334[18:0], v4335[15:0], v5669[19:0]); // 4.0
    wire [31:0] v5670; shift_adder #(18, 30, 1, 1, 32, -13, 0) op_5670 (v4336[17:0], v3256[29:0], v5670[31:0]); // 4.0
    wire [25:0] v5671; shift_adder #(21, 25, 1, 1, 26, -5, 0) op_5671 (v4337[20:0], v2941[24:0], v5671[25:0]); // 4.0
    wire [29:0] v5672; shift_adder #(15, 29, 1, 1, 30, -13, 0) op_5672 (v3308[14:0], v3783[28:0], v5672[29:0]); // 4.0
    wire [28:0] v5673; shift_adder #(28, 25, 1, 1, 29, 2, 0) op_5673 (v2743[27:0], v4338[24:0], v5673[28:0]); // 4.0
    wire [29:0] v5674; shift_adder #(29, 24, 1, 1, 30, 5, 0) op_5674 (v3116[28:0], v4339[23:0], v5674[29:0]); // 4.0
    wire [20:0] v5675; shift_adder #(16, 20, 1, 1, 21, -4, 0) op_5675 (v4340[15:0], v4341[19:0], v5675[20:0]); // 4.0
    wire [38:0] v5676; shift_adder #(37, 20, 1, 1, 39, 18, 0) op_5676 (v4342[36:0], v4343[19:0], v5676[38:0]); // 4.0
    wire [30:0] v5677; shift_adder #(31, 28, 1, 1, 31, 2, 0) op_5677 (v3938[30:0], v3070[27:0], v5677[30:0]); // 4.0
    wire [23:0] v5678; shift_adder #(23, 19, 1, 1, 24, 4, 0) op_5678 (v3168[22:0], v3458[18:0], v5678[23:0]); // 4.0
    wire [17:0] v5679; shift_adder #(17, 14, 1, 1, 18, 2, 0) op_5679 (v3585[16:0], v4344[13:0], v5679[17:0]); // 4.0
    wire [28:0] v5680; shift_adder #(18, 27, 1, 1, 29, -10, 0) op_5680 (v4345[17:0], v4312[26:0], v5680[28:0]); // 4.0
    wire [22:0] v5681; shift_adder #(22, 13, 1, 1, 23, 9, 0) op_5681 (v2997[21:0], v4346[12:0], v5681[22:0]); // 4.0
    wire [28:0] v5682; shift_adder #(22, 28, 1, 1, 29, -7, 0) op_5682 (v4347[21:0], v4348[27:0], v5682[28:0]); // 4.0
    wire [27:0] v5683; shift_adder #(27, 17, 1, 1, 28, 9, 0) op_5683 (v4349[26:0], v3601[16:0], v5683[27:0]); // 4.0
    wire [22:0] v5684; shift_adder #(18, 22, 1, 1, 23, -4, 0) op_5684 (v4350[17:0], v4351[21:0], v5684[22:0]); // 4.0
    wire [20:0] v5685; shift_adder #(18, 21, 1, 1, 21, -2, 0) op_5685 (v3383[17:0], v4352[20:0], v5685[20:0]); // 4.0
    wire [22:0] v5686; shift_adder #(13, 22, 1, 1, 23, -9, 0) op_5686 (v3421[12:0], v4353[21:0], v5686[22:0]); // 4.0
    wire [17:0] v5687; shift_adder #(18, 16, 1, 1, 18, 0, 0) op_5687 (v4354[17:0], v3337[15:0], v5687[17:0]); // 4.0
    wire [18:0] v5688; shift_adder #(16, 18, 1, 1, 19, -1, 0) op_5688 (v4355[15:0], v4356[17:0], v5688[18:0]); // 4.0
    wire [17:0] v5689; shift_adder #(14, 18, 1, 1, 18, -2, 0) op_5689 (v2829[13:0], v4357[17:0], v5689[17:0]); // 4.0
    wire [16:0] v5690; shift_adder #(15, 15, 1, 1, 17, -1, 0) op_5690 (v3666[14:0], v4358[14:0], v5690[16:0]); // 4.0
    wire [15:0] v5691; shift_adder #(14, 14, 1, 1, 16, -1, 0) op_5691 (v4359[13:0], v4360[13:0], v5691[15:0]); // 4.0
    wire [17:0] v5692; shift_adder #(14, 17, 1, 1, 18, -2, 0) op_5692 (v4210[13:0], v4361[16:0], v5692[17:0]); // 4.0
    wire [18:0] v5693; shift_adder #(16, 19, 1, 1, 19, -2, 0) op_5693 (v2977[15:0], v4362[18:0], v5693[18:0]); // 4.0
    wire [21:0] v5694; shift_adder #(18, 20, 1, 1, 22, -3, 0) op_5694 (v3635[17:0], v3777[19:0], v5694[21:0]); // 4.0
    wire [19:0] v5695; shift_adder #(17, 15, 1, 1, 20, 5, 0) op_5695 (v2561[16:0], v4363[14:0], v5695[19:0]); // 4.0
    wire [22:0] v5696; shift_adder #(22, 17, 1, 1, 23, 5, 0) op_5696 (v3007[21:0], v4364[16:0], v5696[22:0]); // 4.0
    wire [24:0] v5697; shift_adder #(14, 23, 1, 1, 25, -10, 0) op_5697 (v4365[13:0], v4366[22:0], v5697[24:0]); // 4.0
    wire [21:0] v5698; shift_adder #(16, 22, 1, 1, 22, -5, 0) op_5698 (v3259[15:0], v4114[21:0], v5698[21:0]); // 4.0
    wire [22:0] v5699; shift_adder #(22, 16, 1, 1, 23, 6, 0) op_5699 (v3036[21:0], v3405[15:0], v5699[22:0]); // 4.0
    wire [24:0] v5700; shift_adder #(23, 24, 1, 1, 25, -2, 0) op_5700 (v4367[22:0], v4058[23:0], v5700[24:0]); // 4.0
    wire [23:0] v5701; shift_adder #(18, 23, 1, 1, 24, -4, 0) op_5701 (v4368[17:0], v3698[22:0], v5701[23:0]); // 4.0
    wire [25:0] v5702; shift_adder #(24, 25, 1, 1, 26, -1, 0) op_5702 (v3807[23:0], v2898[24:0], v5702[25:0]); // 4.0
    wire [31:0] v5703; shift_adder #(23, 30, 1, 1, 32, -8, 0) op_5703 (v4369[22:0], v4370[29:0], v5703[31:0]); // 4.0
    wire [16:0] v5704; shift_adder #(15, 15, 1, 1, 17, 1, 0) op_5704 (v4371[14:0], v4078[14:0], v5704[16:0]); // 4.0
    wire [28:0] v5705; shift_adder #(28, 16, 1, 1, 29, 12, 0) op_5705 (v4372[27:0], v3679[15:0], v5705[28:0]); // 4.0
    wire [24:0] v5706; shift_adder #(23, 25, 1, 1, 25, -1, 0) op_5706 (v4373[22:0], v4164[24:0], v5706[24:0]); // 4.0
    wire [22:0] v5707; shift_adder #(21, 13, 1, 1, 23, 9, 0) op_5707 (v2998[20:0], v4074[12:0], v5707[22:0]); // 4.0
    wire [20:0] v5708; shift_adder #(20, 14, 1, 1, 21, 6, 0) op_5708 (v4374[19:0], v4028[13:0], v5708[20:0]); // 4.0
    wire [27:0] v5709; shift_adder #(26, 16, 1, 1, 28, 11, 0) op_5709 (v4160[25:0], v4375[15:0], v5709[27:0]); // 4.0
    wire [31:0] v5710; shift_adder #(30, 28, 1, 1, 32, 4, 0) op_5710 (v4039[29:0], v3127[27:0], v5710[31:0]); // 4.0
    wire [26:0] v5711; shift_adder #(25, 18, 1, 1, 27, 9, 0) op_5711 (v2959[24:0], v4376[17:0], v5711[26:0]); // 4.0
    wire [33:0] v5712; shift_adder #(13, 18, 1, 1, 34, 16, 1) op_5712 (v4377[12:0], v2474[17:0], v5712[33:0]); // 4.0
    wire [32:0] v5713; shift_adder #(25, 32, 1, 1, 33, -6, 0) op_5713 (v4333[24:0], v3997[31:0], v5713[32:0]); // 4.0
    wire [27:0] v5714; shift_adder #(21, 27, 1, 1, 28, -7, 0) op_5714 (v4378[20:0], v4379[26:0], v5714[27:0]); // 4.0
    wire [39:0] v5715; shift_adder #(31, 39, 1, 1, 40, -8, 0) op_5715 (v3316[30:0], v4380[38:0], v5715[39:0]); // 4.0
    wire [24:0] v5716; shift_adder #(17, 24, 1, 1, 25, -6, 0) op_5716 (v4381[16:0], v4382[23:0], v5716[24:0]); // 4.0
    wire [36:0] v5717; shift_adder #(18, 36, 1, 1, 37, -18, 0) op_5717 (v4269[17:0], v4383[35:0], v5717[36:0]); // 4.0
    wire [37:0] v5718; shift_adder #(37, 17, 1, 1, 38, 21, 0) op_5718 (v4384[36:0], v4385[16:0], v5718[37:0]); // 4.0
    wire [14:0] v5719; shift_adder #(14, 13, 1, 1, 15, 0, 0) op_5719 (v3096[13:0], v4386[12:0], v5719[14:0]); // 4.0
    wire [27:0] v5720; shift_adder #(27, 17, 1, 1, 28, 9, 0) op_5720 (v2538[26:0], v4387[16:0], v5720[27:0]); // 4.0
    wire [30:0] v5721; shift_adder #(31, 19, 1, 1, 31, 10, 0) op_5721 (v4388[30:0], v3376[18:0], v5721[30:0]); // 4.0
    wire [20:0] v5722; shift_adder #(19, 17, 1, 1, 21, 3, 0) op_5722 (v4389[18:0], v3288[16:0], v5722[20:0]); // 4.0
    wire [25:0] v5723; shift_adder #(26, 17, 1, 1, 26, 6, 0) op_5723 (v4390[25:0], v4391[16:0], v5723[25:0]); // 4.0
    wire [27:0] v5724; shift_adder #(17, 25, 1, 1, 28, -11, 0) op_5724 (v4392[16:0], v4393[24:0], v5724[27:0]); // 4.0
    wire [20:0] v5725; shift_adder #(16, 19, 1, 1, 21, -5, 0) op_5725 (v2614[15:0], v4007[18:0], v5725[20:0]); // 4.0
    wire [21:0] v5726; shift_adder #(20, 21, 1, 1, 22, -1, 0) op_5726 (v4394[19:0], v4395[20:0], v5726[21:0]); // 4.0
    wire [24:0] v5727; shift_adder #(25, 14, 1, 1, 25, 9, 0) op_5727 (v4396[24:0], v2848[13:0], v5727[24:0]); // 4.0
    wire [17:0] v5728; shift_adder #(15, 17, 1, 1, 18, -2, 0) op_5728 (v3696[14:0], v3274[16:0], v5728[17:0]); // 4.0
    wire [18:0] v5729; shift_adder #(17, 17, 1, 1, 19, -1, 0) op_5729 (v4397[16:0], v4293[16:0], v5729[18:0]); // 4.0
    wire [21:0] v5730; shift_adder #(21, 20, 1, 1, 22, 1, 0) op_5730 (v4398[20:0], v4399[19:0], v5730[21:0]); // 4.0
    wire [16:0] v5731; shift_adder #(14, 15, 1, 1, 17, -3, 0) op_5731 (v4400[13:0], v4401[14:0], v5731[16:0]); // 4.0
    wire [23:0] v5732; shift_adder #(19, 23, 1, 1, 24, -4, 0) op_5732 (v2544[18:0], v4402[22:0], v5732[23:0]); // 4.0
    wire [29:0] v5733; shift_adder #(27, 24, 1, 1, 30, 6, 0) op_5733 (v4403[26:0], v4404[23:0], v5733[29:0]); // 4.0
    wire [28:0] v5734; shift_adder #(27, 28, 1, 1, 29, 0, 0) op_5734 (v4405[26:0], v4406[27:0], v5734[28:0]); // 4.0
    wire [24:0] v5735; shift_adder #(23, 18, 1, 1, 25, 6, 0) op_5735 (v4407[22:0], v4350[17:0], v5735[24:0]); // 4.0
    wire [25:0] v5736; shift_adder #(25, 20, 1, 1, 26, 6, 0) op_5736 (v3517[24:0], v4408[19:0], v5736[25:0]); // 4.0
    wire [21:0] v5737; shift_adder #(18, 21, 1, 1, 22, -3, 0) op_5737 (v4409[17:0], v2746[20:0], v5737[21:0]); // 4.0
    wire [17:0] v5738; shift_adder #(14, 18, 1, 1, 18, -2, 0) op_5738 (v3923[13:0], v4410[17:0], v5738[17:0]); // 4.0
    wire [14:0] v5739; shift_adder #(14, 15, 1, 1, 15, 0, 0) op_5739 (v3252[13:0], v4411[14:0], v5739[14:0]); // 4.0
    wire [22:0] v5740; shift_adder #(21, 22, 1, 1, 23, -1, 0) op_5740 (v3731[20:0], v4412[21:0], v5740[22:0]); // 4.0
    wire [29:0] v5741; shift_adder #(29, 18, 1, 1, 30, 12, 0) op_5741 (v4413[28:0], v3719[17:0], v5741[29:0]); // 4.0
    wire [22:0] v5742; shift_adder #(16, 22, 1, 1, 23, -6, 0) op_5742 (v2863[15:0], v4414[21:0], v5742[22:0]); // 4.0
    wire [29:0] v5743; shift_adder #(28, 29, 1, 1, 30, -1, 0) op_5743 (v4415[27:0], v2946[28:0], v5743[29:0]); // 4.0
    wire [32:0] v5744; shift_adder #(32, 29, 1, 1, 33, 4, 0) op_5744 (v2742[31:0], v3579[28:0], v5744[32:0]); // 4.0
    wire [36:0] v5745; shift_adder #(36, 24, 1, 1, 37, 12, 0) op_5745 (v4416[35:0], v4417[23:0], v5745[36:0]); // 4.0
    wire [16:0] v5746; shift_adder #(16, 15, 1, 1, 17, 0, 0) op_5746 (v4418[15:0], v4419[14:0], v5746[16:0]); // 4.0
    wire [17:0] v5747; shift_adder #(13, 17, 1, 1, 18, -2, 0) op_5747 (v4420[12:0], v4421[16:0], v5747[17:0]); // 4.0
    wire [19:0] v5748; shift_adder #(17, 18, 1, 1, 20, -2, 0) op_5748 (v4133[16:0], v4422[17:0], v5748[19:0]); // 4.0
    wire [21:0] v5749; shift_adder #(21, 15, 1, 1, 22, 6, 0) op_5749 (v2592[20:0], v4423[14:0], v5749[21:0]); // 4.0
    wire [16:0] v5750; shift_adder #(16, 15, 1, 1, 17, 1, 0) op_5750 (v3621[15:0], v4424[14:0], v5750[16:0]); // 4.0
    wire [17:0] v5751; shift_adder #(14, 17, 1, 1, 18, -1, 0) op_5751 (v4425[13:0], v4426[16:0], v5751[17:0]); // 4.0
    wire [19:0] v5752; shift_adder #(16, 19, 1, 1, 20, -3, 0) op_5752 (v3596[15:0], v4428[18:0], v5752[19:0]); // 4.0
    wire [27:0] v5753; shift_adder #(15, 27, 1, 1, 28, -11, 0) op_5753 (v3582[14:0], v4379[26:0], v5753[27:0]); // 4.0
    wire [36:0] v5754; shift_adder #(14, 12, 1, 1, 37, 25, 1) op_5754 (v4177[13:0], v2502[11:0], v5754[36:0]); // 4.0
    wire [35:0] v5755; shift_adder #(35, 20, 1, 1, 36, 15, 0) op_5755 (v4429[34:0], v4430[19:0], v5755[35:0]); // 4.0
    wire [33:0] v5756; shift_adder #(34, 14, 1, 1, 34, 18, 0) op_5756 (v4431[33:0], v2526[13:0], v5756[33:0]); // 4.0
    wire [37:0] v5757; shift_adder #(26, 35, 1, 1, 38, -12, 0) op_5757 (v3004[25:0], v3788[34:0], v5757[37:0]); // 4.0
    wire [31:0] v5758; shift_adder #(31, 22, 1, 1, 32, 8, 0) op_5758 (v4432[30:0], v3072[21:0], v5758[31:0]); // 4.0
    wire [25:0] v5759; shift_adder #(26, 13, 1, 1, 26, 11, 0) op_5759 (v4168[25:0], v4433[12:0], v5759[25:0]); // 4.0
    wire [24:0] v5760; shift_adder #(23, 24, 1, 1, 25, -2, 0) op_5760 (v4434[22:0], v3824[23:0], v5760[24:0]); // 4.0
    wire [18:0] v5761; shift_adder #(18, 16, 1, 1, 19, 1, 0) op_5761 (v2611[17:0], v4435[15:0], v5761[18:0]); // 4.0
    wire [27:0] v5762; shift_adder #(24, 26, 1, 1, 28, -3, 0) op_5762 (v4436[23:0], v3983[25:0], v5762[27:0]); // 4.0
    wire [25:0] v5763; shift_adder #(24, 26, 1, 1, 26, 0, 0) op_5763 (v4437[23:0], v4438[25:0], v5763[25:0]); // 4.0
    wire [31:0] v5764; shift_adder #(20, 30, 1, 1, 32, -12, 0) op_5764 (v3158[19:0], v4439[29:0], v5764[31:0]); // 4.0
    wire [14:0] v5765; shift_adder #(13, 14, 1, 1, 15, -1, 0) op_5765 (v4440[12:0], v3369[13:0], v5765[14:0]); // 4.0
    wire [29:0] v5766; shift_adder #(30, 17, 1, 1, 30, 11, 0) op_5766 (v3348[29:0], v3733[16:0], v5766[29:0]); // 4.0
    wire [24:0] v5767; shift_adder #(24, 24, 1, 1, 25, 0, 0) op_5767 (v4035[23:0], v3510[23:0], v5767[24:0]); // 4.0
    wire [16:0] v5768; shift_adder #(17, 15, 1, 1, 17, 1, 0) op_5768 (v4441[16:0], v4442[14:0], v5768[16:0]); // 4.0
    wire [19:0] v5769; shift_adder #(20, 14, 1, 1, 20, 3, 0) op_5769 (v4443[19:0], v4187[13:0], v5769[19:0]); // 4.0
    wire [19:0] v5770; shift_adder #(16, 18, 1, 1, 20, -4, 0) op_5770 (v4444[15:0], v3928[17:0], v5770[19:0]); // 4.0
    wire [24:0] v5771; shift_adder #(21, 25, 1, 1, 25, -2, 0) op_5771 (v4445[20:0], v4446[24:0], v5771[24:0]); // 5.0
    wire [24:0] v5772; shift_adder #(23, 25, 1, 1, 25, -1, 0) op_5772 (v4447[22:0], v4448[24:0], v5772[24:0]); // 5.0
    wire [25:0] v5773; shift_adder #(11, 26, 1, 1, 26, -3, 1) op_5773 (v152[10:0], v4449[25:0], v5773[25:0]); // 5.0
    wire [29:0] v5774; shift_adder #(27, 25, 1, 1, 30, 4, 0) op_5774 (v4450[26:0], v4451[24:0], v5774[29:0]); // 5.0
    wire [32:0] v5775; shift_adder #(9, 28, 1, 1, 33, -23, 1) op_5775 (v128[8:0], v4452[27:0], v5775[32:0]); // 5.0
    wire [25:0] v5776; shift_adder #(25, 18, 1, 1, 26, 7, 0) op_5776 (v4453[24:0], v4454[17:0], v5776[25:0]); // 5.0
    wire [31:0] v5777; shift_adder #(28, 31, 1, 1, 32, 0, 0) op_5777 (v4455[27:0], v4456[30:0], v5777[31:0]); // 5.0
    wire [26:0] v5778; shift_adder #(27, 17, 1, 1, 27, 8, 0) op_5778 (v4457[26:0], v4458[16:0], v5778[26:0]); // 5.0
    wire [28:0] v5779; shift_adder #(23, 28, 1, 1, 29, -6, 0) op_5779 (v4459[22:0], v4460[27:0], v5779[28:0]); // 5.0
    wire [32:0] v5780; shift_adder #(32, 19, 1, 1, 33, 12, 0) op_5780 (v4461[31:0], v4462[18:0], v5780[32:0]); // 5.0
    wire [25:0] v5781; shift_adder #(22, 25, 1, 1, 26, -4, 0) op_5781 (v4463[21:0], v4464[24:0], v5781[25:0]); // 5.0
    wire [18:0] v5782; shift_adder #(15, 16, 1, 1, 19, 3, 0) op_5782 (v4465[14:0], v4466[15:0], v5782[18:0]); // 5.0
    wire [24:0] v5783; shift_adder #(24, 20, 1, 1, 25, 4, 0) op_5783 (v4468[23:0], v4469[19:0], v5783[24:0]); // 5.0
    wire [29:0] v5784; shift_adder #(27, 29, 1, 1, 30, -1, 0) op_5784 (v4470[26:0], v4471[28:0], v5784[29:0]); // 5.0
    wire [23:0] v5785; shift_adder #(21, 23, 1, 1, 24, -2, 0) op_5785 (v4472[20:0], v4473[22:0], v5785[23:0]); // 5.0
    wire [22:0] v5786; shift_adder #(22, 18, 1, 1, 23, 4, 0) op_5786 (v4474[21:0], v4475[17:0], v5786[22:0]); // 5.0
    wire [31:0] v5787; shift_adder #(31, 29, 1, 1, 32, 0, 0) op_5787 (v4476[30:0], v4477[28:0], v5787[31:0]); // 5.0
    wire [36:0] v5788; shift_adder #(35, 17, 1, 1, 37, -2, 1) op_5788 (v4478[34:0], v4479[16:0], v5788[36:0]); // 5.0
    wire [32:0] v5789; shift_adder #(15, 32, 1, 1, 33, -17, 0) op_5789 (v4480[14:0], v4481[31:0], v5789[32:0]); // 5.0
    wire [22:0] v5790; shift_adder #(23, 20, 1, 1, 23, 2, 0) op_5790 (v4482[22:0], v4483[19:0], v5790[22:0]); // 5.0
    wire [19:0] v5791; shift_adder #(19, 19, 1, 1, 20, 1, 0) op_5791 (v4484[18:0], v4485[18:0], v5791[19:0]); // 5.0
    wire [31:0] v5792; shift_adder #(8, 19, 1, 1, 32, 13, 1) op_5792 (v125[7:0], v4486[18:0], v5792[31:0]); // 5.0
    wire [26:0] v5793; shift_adder #(22, 25, 1, 1, 27, -5, 0) op_5793 (v4487[21:0], v4488[24:0], v5793[26:0]); // 5.0
    wire [22:0] v5794; shift_adder #(21, 22, 1, 1, 23, -2, 0) op_5794 (v4489[20:0], v4490[21:0], v5794[22:0]); // 5.0
    wire [22:0] v5795; shift_adder #(22, 16, 1, 1, 23, 6, 0) op_5795 (v4491[21:0], v4492[15:0], v5795[22:0]); // 5.0
    wire [20:0] v5796; shift_adder #(17, 20, 1, 1, 21, -2, 0) op_5796 (v4493[16:0], v4494[19:0], v5796[20:0]); // 5.0
    wire [25:0] v5797; shift_adder #(20, 20, 1, 1, 26, 5, 0) op_5797 (v4495[19:0], v4496[19:0], v5797[25:0]); // 5.0
    wire [26:0] v5798; shift_adder #(21, 27, 1, 1, 27, -2, 0) op_5798 (v4497[20:0], v4498[26:0], v5798[26:0]); // 5.0
    wire [29:0] v5799; shift_adder #(23, 29, 1, 1, 30, -5, 0) op_5799 (v4499[22:0], v4500[28:0], v5799[29:0]); // 5.0
    wire [34:0] v5800; shift_adder #(11, 35, 1, 1, 35, -5, 1) op_5800 (v185[10:0], v4501[34:0], v5800[34:0]); // 5.0
    wire [23:0] v5801; shift_adder #(23, 20, 1, 1, 24, 3, 0) op_5801 (v4502[22:0], v4503[19:0], v5801[23:0]); // 5.0
    wire [17:0] v5802; shift_adder #(8, 17, 1, 1, 18, -7, 1) op_5802 (v69[7:0], v4504[16:0], v5802[17:0]); // 5.0
    wire [27:0] v5803; shift_adder #(23, 26, 1, 1, 28, -4, 0) op_5803 (v4505[22:0], v4506[25:0], v5803[27:0]); // 5.0
    wire [27:0] v5804; shift_adder #(20, 27, 1, 1, 28, -6, 0) op_5804 (v4507[19:0], v4508[26:0], v5804[27:0]); // 5.0
    wire [29:0] v5805; shift_adder #(20, 28, 1, 1, 30, -10, 0) op_5805 (v4509[19:0], v4510[27:0], v5805[29:0]); // 5.0
    wire [32:0] v5806; shift_adder #(31, 20, 1, 1, 33, 13, 0) op_5806 (v4511[30:0], v4512[19:0], v5806[32:0]); // 5.0
    wire [34:0] v5807; shift_adder #(23, 34, 1, 1, 35, -10, 0) op_5807 (v4513[22:0], v4514[33:0], v5807[34:0]); // 5.0
    wire [28:0] v5808; shift_adder #(28, 26, 1, 1, 29, 2, 0) op_5808 (v4515[27:0], v4516[25:0], v5808[28:0]); // 5.0
    wire [36:0] v5809; shift_adder #(36, 17, 1, 1, 37, -1, 1) op_5809 (v4517[35:0], v4518[16:0], v5809[36:0]); // 5.0
    wire [19:0] v5810; shift_adder #(18, 18, 1, 1, 20, -1, 0) op_5810 (v4519[17:0], v4520[17:0], v5810[19:0]); // 5.0
    wire [23:0] v5811; shift_adder #(19, 22, 1, 1, 24, -4, 0) op_5811 (v4521[18:0], v4522[21:0], v5811[23:0]); // 5.0
    wire [21:0] v5812; shift_adder #(21, 19, 1, 1, 22, 0, 0) op_5812 (v4523[20:0], v4524[18:0], v5812[21:0]); // 5.0
    wire [19:0] v5813; shift_adder #(16, 20, 1, 1, 20, -2, 0) op_5813 (v4525[15:0], v4526[19:0], v5813[19:0]); // 5.0
    wire [27:0] v5814; shift_adder #(27, 20, 1, 1, 28, 7, 0) op_5814 (v4528[26:0], v4529[19:0], v5814[27:0]); // 5.0
    wire [39:0] v5815; shift_adder #(39, 38, 1, 1, 40, 1, 0) op_5815 (v4530[38:0], v4531[37:0], v5815[39:0]); // 5.0
    wire [28:0] v5816; shift_adder #(28, 15, 1, 1, 29, 13, 0) op_5816 (v4532[27:0], v4533[14:0], v5816[28:0]); // 5.0
    wire [24:0] v5817; shift_adder #(24, 23, 1, 1, 25, 0, 0) op_5817 (v4534[23:0], v4535[22:0], v5817[24:0]); // 5.0
    wire [24:0] v5818; shift_adder #(24, 23, 1, 1, 25, -1, 0) op_5818 (v4536[23:0], v4537[22:0], v5818[24:0]); // 5.0
    wire [24:0] v5819; shift_adder #(25, 14, 1, 1, 25, 9, 0) op_5819 (v4538[24:0], v4539[13:0], v5819[24:0]); // 5.0
    wire [26:0] v5820; shift_adder #(25, 23, 1, 1, 27, 3, 0) op_5820 (v4540[24:0], v4541[22:0], v5820[26:0]); // 5.0
    wire [30:0] v5821; shift_adder #(26, 30, 1, 1, 31, -3, 0) op_5821 (v4542[25:0], v4543[29:0], v5821[30:0]); // 5.0
    wire [28:0] v5822; shift_adder #(27, 23, 1, 1, 29, 5, 0) op_5822 (v4544[26:0], v4545[22:0], v5822[28:0]); // 5.0
    wire [25:0] v5823; shift_adder #(26, 17, 1, 1, 26, 8, 0) op_5823 (v4546[25:0], v4547[16:0], v5823[25:0]); // 5.0
    wire [36:0] v5824; shift_adder #(35, 31, 1, 1, 37, 5, 0) op_5824 (v4548[34:0], v4549[30:0], v5824[36:0]); // 5.0
    wire [27:0] v5825; shift_adder #(20, 27, 1, 1, 28, -8, 0) op_5825 (v4550[19:0], v4551[26:0], v5825[27:0]); // 5.0
    wire [23:0] v5826; shift_adder #(23, 21, 1, 1, 24, 2, 0) op_5826 (v4552[22:0], v4553[20:0], v5826[23:0]); // 5.0
    wire [23:0] v5827; shift_adder #(20, 23, 1, 1, 24, -3, 0) op_5827 (v4554[19:0], v4555[22:0], v5827[23:0]); // 5.0
    wire [31:0] v5828; shift_adder #(8, 32, 1, 1, 32, -19, 1) op_5828 (v102[7:0], v4556[31:0], v5828[31:0]); // 5.0
    wire [27:0] v5829; shift_adder #(28, 17, 1, 1, 28, 8, 0) op_5829 (v4557[27:0], v4558[16:0], v5829[27:0]); // 5.0
    wire [40:0] v5830; shift_adder #(39, 35, 1, 1, 41, 5, 0) op_5830 (v4559[38:0], v4560[34:0], v5830[40:0]); // 5.0
    wire [18:0] v5831; shift_adder #(17, 17, 1, 1, 19, -2, 0) op_5831 (v4561[16:0], v4562[16:0], v5831[18:0]); // 5.0
    wire [34:0] v5832; shift_adder #(32, 34, 1, 1, 35, -3, 0) op_5832 (v4563[31:0], v4564[33:0], v5832[34:0]); // 5.0
    wire [36:0] v5833; shift_adder #(26, 37, 1, 1, 37, -10, 0) op_5833 (v4565[25:0], v4566[36:0], v5833[36:0]); // 5.0
    wire [23:0] v5834; shift_adder #(23, 17, 1, 1, 24, 5, 0) op_5834 (v4567[22:0], v4568[16:0], v5834[23:0]); // 5.0
    wire [29:0] v5835; shift_adder #(21, 28, 1, 1, 30, -8, 0) op_5835 (v4569[20:0], v4570[27:0], v5835[29:0]); // 5.0
    wire [20:0] v5836; shift_adder #(19, 19, 1, 1, 21, -2, 0) op_5836 (v4571[18:0], v4572[18:0], v5836[20:0]); // 5.0
    wire [18:0] v5837; shift_adder #(19, 16, 1, 1, 19, 0, 0) op_5837 (v4573[18:0], v4574[15:0], v5837[18:0]); // 5.0
    wire [28:0] v5838; shift_adder #(27, 22, 1, 1, 29, 6, 0) op_5838 (v4575[26:0], v4576[21:0], v5838[28:0]); // 5.0
    wire [32:0] v5839; shift_adder #(29, 31, 1, 1, 33, -3, 0) op_5839 (v4577[28:0], v4578[30:0], v5839[32:0]); // 5.0
    wire [33:0] v5840; shift_adder #(27, 33, 1, 1, 34, -6, 0) op_5840 (v4579[26:0], v4580[32:0], v5840[33:0]); // 5.0
    wire [28:0] v5841; shift_adder #(27, 29, 1, 1, 29, 0, 0) op_5841 (v4470[26:0], v4581[28:0], v5841[28:0]); // 5.0
    wire [23:0] v5842; shift_adder #(22, 17, 1, 1, 24, 7, 0) op_5842 (v4582[21:0], v4583[16:0], v5842[23:0]); // 5.0
    wire [22:0] v5843; shift_adder #(20, 22, 1, 1, 23, 1, 0) op_5843 (v4584[19:0], v4585[21:0], v5843[22:0]); // 5.0
    wire [37:0] v5844; shift_adder #(37, 27, 1, 1, 38, 9, 0) op_5844 (v4586[36:0], v4587[26:0], v5844[37:0]); // 5.0
    wire [19:0] v5845; shift_adder #(17, 20, 1, 1, 20, -1, 0) op_5845 (v4588[16:0], v4589[19:0], v5845[19:0]); // 5.0
    wire [19:0] v5846; shift_adder #(19, 18, 1, 1, 20, 1, 0) op_5846 (v4590[18:0], v4591[17:0], v5846[19:0]); // 5.0
    wire [21:0] v5847; shift_adder #(18, 21, 1, 1, 22, -1, 0) op_5847 (v4592[17:0], v4593[20:0], v5847[21:0]); // 5.0
    wire [25:0] v5848; shift_adder #(23, 25, 1, 1, 26, 1, 0) op_5848 (v4594[22:0], v4595[24:0], v5848[25:0]); // 5.0
    wire [33:0] v5849; shift_adder #(33, 20, 1, 1, 34, 13, 0) op_5849 (v4596[32:0], v4597[19:0], v5849[33:0]); // 5.0
    wire [31:0] v5850; shift_adder #(31, 26, 1, 1, 32, 4, 0) op_5850 (v4598[30:0], v4599[25:0], v5850[31:0]); // 5.0
    wire [31:0] v5851; shift_adder #(25, 31, 1, 1, 32, -5, 0) op_5851 (v4600[24:0], v4601[30:0], v5851[31:0]); // 5.0
    wire [27:0] v5852; shift_adder #(25, 27, 1, 1, 28, -2, 0) op_5852 (v4602[24:0], v4603[26:0], v5852[27:0]); // 5.0
    wire [19:0] v5853; shift_adder #(13, 20, 1, 1, 20, -6, 1) op_5853 (v346[12:0], v4604[19:0], v5853[19:0]); // 5.0
    wire [29:0] v5854; shift_adder #(17, 30, 1, 1, 30, -12, 0) op_5854 (v4605[16:0], v4606[29:0], v5854[29:0]); // 5.0
    wire [37:0] v5855; shift_adder #(38, 17, 1, 1, 38, 0, 1) op_5855 (v4607[37:0], v4608[16:0], v5855[37:0]); // 5.0
    wire [19:0] v5856; shift_adder #(18, 19, 1, 1, 20, 0, 0) op_5856 (v4609[17:0], v4610[18:0], v5856[19:0]); // 5.0
    wire [32:0] v5857; shift_adder #(29, 32, 1, 1, 33, -2, 0) op_5857 (v4611[28:0], v4612[31:0], v5857[32:0]); // 5.0
    wire [29:0] v5858; shift_adder #(29, 26, 1, 1, 30, 3, 0) op_5858 (v4613[28:0], v4614[25:0], v5858[29:0]); // 5.0
    wire [23:0] v5859; shift_adder #(23, 18, 1, 1, 24, 5, 0) op_5859 (v4552[22:0], v4615[17:0], v5859[23:0]); // 5.0
    wire [23:0] v5860; shift_adder #(22, 22, 1, 1, 24, -2, 0) op_5860 (v4616[21:0], v4617[21:0], v5860[23:0]); // 5.0
    wire [32:0] v5861; shift_adder #(17, 31, 1, 1, 33, -15, 0) op_5861 (v4618[16:0], v4511[30:0], v5861[32:0]); // 5.0
    wire [36:0] v5862; shift_adder #(33, 36, 1, 1, 37, -3, 0) op_5862 (v4619[32:0], v4620[35:0], v5862[36:0]); // 5.0
    wire [37:0] v5863; shift_adder #(36, 33, 1, 1, 38, 4, 0) op_5863 (v4621[35:0], v4622[32:0], v5863[37:0]); // 5.0
    wire [30:0] v5864; shift_adder #(18, 30, 1, 1, 31, -11, 0) op_5864 (v4623[17:0], v4624[29:0], v5864[30:0]); // 5.0
    wire [32:0] v5865; shift_adder #(27, 31, 1, 1, 33, -5, 0) op_5865 (v4551[26:0], v4625[30:0], v5865[32:0]); // 5.0
    wire [31:0] v5866; shift_adder #(31, 26, 1, 1, 32, 5, 0) op_5866 (v4626[30:0], v4627[25:0], v5866[31:0]); // 5.0
    wire [23:0] v5867; shift_adder #(23, 21, 1, 1, 24, 3, 0) op_5867 (v4628[22:0], v4629[20:0], v5867[23:0]); // 5.0
    wire [30:0] v5868; shift_adder #(25, 30, 1, 1, 31, -6, 0) op_5868 (v4630[24:0], v4631[29:0], v5868[30:0]); // 5.0
    wire [21:0] v5869; shift_adder #(20, 20, 1, 1, 22, 1, 0) op_5869 (v4632[19:0], v4633[19:0], v5869[21:0]); // 5.0
    wire [27:0] v5870; shift_adder #(24, 28, 1, 1, 28, -2, 0) op_5870 (v4634[23:0], v4635[27:0], v5870[27:0]); // 5.0
    wire [30:0] v5871; shift_adder #(30, 22, 1, 1, 31, 8, 0) op_5871 (v4636[29:0], v4637[21:0], v5871[30:0]); // 5.0
    wire [33:0] v5872; shift_adder #(32, 23, 1, 1, 34, 11, 0) op_5872 (v4638[31:0], v4639[22:0], v5872[33:0]); // 5.0
    wire [18:0] v5873; shift_adder #(15, 19, 1, 1, 19, -1, 0) op_5873 (v4640[14:0], v4641[18:0], v5873[18:0]); // 5.0
    wire [31:0] v5874; shift_adder #(31, 26, 1, 1, 32, 6, 0) op_5874 (v4643[30:0], v4644[25:0], v5874[31:0]); // 5.0
    wire [26:0] v5875; shift_adder #(24, 27, 1, 1, 27, -2, 0) op_5875 (v4645[23:0], v4544[26:0], v5875[26:0]); // 5.0
    wire [32:0] v5876; shift_adder #(31, 32, 1, 1, 33, -1, 0) op_5876 (v4646[30:0], v4647[31:0], v5876[32:0]); // 5.0
    wire [35:0] v5877; shift_adder #(17, 29, 1, 1, 36, 7, 1) op_5877 (v4648[16:0], v2861[28:0], v5877[35:0]); // 5.0
    wire [33:0] v5878; shift_adder #(33, 19, 1, 1, 34, 15, 0) op_5878 (v4649[32:0], v4650[18:0], v5878[33:0]); // 5.0
    wire [30:0] v5879; shift_adder #(30, 26, 1, 1, 31, 4, 0) op_5879 (v4651[29:0], v4652[25:0], v5879[30:0]); // 5.0
    wire [34:0] v5880; shift_adder #(34, 19, 1, 1, 35, 15, 0) op_5880 (v4653[33:0], v4654[18:0], v5880[34:0]); // 5.0
    wire [20:0] v5881; shift_adder #(17, 19, 1, 1, 21, -3, 0) op_5881 (v4655[16:0], v4656[18:0], v5881[20:0]); // 5.0
    wire [35:0] v5882; shift_adder #(35, 17, 1, 1, 36, -1, 1) op_5882 (v4657[34:0], v4658[16:0], v5882[35:0]); // 5.0
    wire [40:0] v5883; shift_adder #(40, 29, 1, 1, 41, 10, 0) op_5883 (v4659[39:0], v4660[28:0], v5883[40:0]); // 5.0
    wire [28:0] v5884; shift_adder #(26, 28, 1, 1, 29, -3, 0) op_5884 (v4661[25:0], v4662[27:0], v5884[28:0]); // 5.0
    wire [32:0] v5885; shift_adder #(31, 24, 1, 1, 33, 9, 0) op_5885 (v4663[30:0], v4664[23:0], v5885[32:0]); // 5.0
    wire [28:0] v5886; shift_adder #(22, 29, 1, 1, 29, -5, 0) op_5886 (v4665[21:0], v4666[28:0], v5886[28:0]); // 5.0
    wire [31:0] v5887; shift_adder #(32, 30, 1, 1, 32, 0, 0) op_5887 (v4667[31:0], v4668[29:0], v5887[31:0]); // 5.0
    wire [17:0] v5888; shift_adder #(16, 17, 1, 1, 18, -1, 0) op_5888 (v4669[15:0], v4670[16:0], v5888[17:0]); // 5.0
    wire [24:0] v5889; shift_adder #(24, 21, 1, 1, 25, 2, 0) op_5889 (v4671[23:0], v4672[20:0], v5889[24:0]); // 5.0
    wire [25:0] v5890; shift_adder #(25, 23, 1, 1, 26, 1, 0) op_5890 (v4673[24:0], v4674[22:0], v5890[25:0]); // 5.0
    wire [21:0] v5891; shift_adder #(22, 18, 1, 1, 22, 1, 0) op_5891 (v4675[21:0], v4676[17:0], v5891[21:0]); // 5.0
    wire [28:0] v5892; shift_adder #(26, 16, 1, 1, 29, 12, 0) op_5892 (v4677[25:0], v4678[15:0], v5892[28:0]); // 5.0
    wire [24:0] v5893; shift_adder #(21, 21, 1, 1, 25, 4, 0) op_5893 (v4679[20:0], v4680[20:0], v5893[24:0]); // 5.0
    wire [24:0] v5894; shift_adder #(23, 24, 1, 1, 25, -1, 0) op_5894 (v4681[22:0], v4682[23:0], v5894[24:0]); // 5.0
    wire [19:0] v5895; shift_adder #(19, 16, 1, 1, 20, 2, 0) op_5895 (v4610[18:0], v4492[15:0], v5895[19:0]); // 5.0
    wire [20:0] v5896; shift_adder #(20, 20, 1, 1, 21, 0, 0) op_5896 (v4683[19:0], v4684[19:0], v5896[20:0]); // 5.0
    wire [20:0] v5897; shift_adder #(20, 19, 1, 1, 21, 0, 0) op_5897 (v4685[19:0], v4686[18:0], v5897[20:0]); // 5.0
    wire [32:0] v5898; shift_adder #(33, 29, 1, 1, 33, 2, 0) op_5898 (v4687[32:0], v4688[28:0], v5898[32:0]); // 5.0
    wire [34:0] v5899; shift_adder #(29, 34, 1, 1, 35, -6, 0) op_5899 (v4689[28:0], v4690[33:0], v5899[34:0]); // 5.0
    wire [32:0] v5900; shift_adder #(33, 24, 1, 1, 33, 6, 0) op_5900 (v4691[32:0], v4692[23:0], v5900[32:0]); // 5.0
    wire [22:0] v5901; shift_adder #(20, 22, 1, 1, 23, -2, 0) op_5901 (v4693[19:0], v4637[21:0], v5901[22:0]); // 5.0
    wire [17:0] v5902; shift_adder #(16, 17, 1, 1, 18, -1, 0) op_5902 (v4694[15:0], v4695[16:0], v5902[17:0]); // 5.0
    wire [23:0] v5903; shift_adder #(17, 24, 1, 1, 24, -5, 0) op_5903 (v4697[16:0], v4698[23:0], v5903[23:0]); // 5.0
    wire [36:0] v5904; shift_adder #(35, 27, 1, 1, 37, 9, 0) op_5904 (v4699[34:0], v4700[26:0], v5904[36:0]); // 5.0
    wire [32:0] v5905; shift_adder #(25, 30, 1, 1, 33, -7, 0) op_5905 (v4701[24:0], v4702[29:0], v5905[32:0]); // 5.0
    wire [26:0] v5906; shift_adder #(21, 24, 1, 1, 27, -5, 0) op_5906 (v4703[20:0], v4704[23:0], v5906[26:0]); // 5.0
    wire [23:0] v5907; shift_adder #(24, 15, 1, 1, 24, 6, 0) op_5907 (v4705[23:0], v4706[14:0], v5907[23:0]); // 5.0
    wire [20:0] v5908; shift_adder #(21, 18, 1, 1, 21, 2, 0) op_5908 (v4707[20:0], v4708[17:0], v5908[20:0]); // 5.0
    wire [31:0] v5909; shift_adder #(31, 15, 1, 1, 32, 17, 0) op_5909 (v4709[30:0], v4710[14:0], v5909[31:0]); // 5.0
    wire [19:0] v5910; shift_adder #(11, 19, 1, 1, 20, -9, 0) op_5910 (v294[10:0], v4711[18:0], v5910[19:0]); // 5.0
    wire [30:0] v5911; shift_adder #(26, 30, 1, 1, 31, -3, 0) op_5911 (v4712[25:0], v4713[29:0], v5911[30:0]); // 5.0
    wire [33:0] v5912; shift_adder #(8, 32, 1, 1, 34, 2, 0) op_5912 (v114[7:0], v4714[31:0], v5912[33:0]); // 5.0
    wire [38:0] v5913; shift_adder #(17, 17, 1, 1, 39, 22, 1) op_5913 (v4715[16:0], v2968[16:0], v5913[38:0]); // 5.0
    wire [41:0] v5914; shift_adder #(39, 41, 1, 1, 42, -2, 0) op_5914 (v4716[38:0], v4717[40:0], v5914[41:0]); // 5.0
    wire [19:0] v5915; shift_adder #(19, 15, 1, 1, 20, 1, 0) op_5915 (v4718[18:0], v4719[14:0], v5915[19:0]); // 5.0
    wire [18:0] v5916; shift_adder #(17, 17, 1, 1, 19, -1, 0) op_5916 (v4720[16:0], v4721[16:0], v5916[18:0]); // 5.0
    wire [22:0] v5917; shift_adder #(17, 23, 1, 1, 23, -3, 0) op_5917 (v4722[16:0], v4723[22:0], v5917[22:0]); // 5.0
    wire [21:0] v5918; shift_adder #(20, 16, 1, 1, 22, 6, 0) op_5918 (v4724[19:0], v4725[15:0], v5918[21:0]); // 5.0
    wire [21:0] v5919; shift_adder #(22, 18, 1, 1, 22, 3, 0) op_5919 (v4726[21:0], v4727[17:0], v5919[21:0]); // 5.0
    wire [26:0] v5920; shift_adder #(26, 20, 1, 1, 27, 5, 0) op_5920 (v4728[25:0], v4729[19:0], v5920[26:0]); // 5.0
    wire [25:0] v5921; shift_adder #(17, 26, 1, 1, 26, -7, 0) op_5921 (v4730[16:0], v4731[25:0], v5921[25:0]); // 5.0
    wire [24:0] v5922; shift_adder #(22, 23, 1, 1, 25, 2, 0) op_5922 (v4732[21:0], v4733[22:0], v5922[24:0]); // 5.0
    wire [24:0] v5923; shift_adder #(24, 23, 1, 1, 25, 1, 0) op_5923 (v4734[23:0], v4735[22:0], v5923[24:0]); // 5.0
    wire [33:0] v5924; shift_adder #(31, 28, 1, 1, 34, 6, 0) op_5924 (v4736[30:0], v4737[27:0], v5924[33:0]); // 5.0
    wire [36:0] v5925; shift_adder #(23, 36, 1, 1, 37, -13, 0) op_5925 (v4738[22:0], v4739[35:0], v5925[36:0]); // 5.0
    wire [22:0] v5926; shift_adder #(23, 18, 1, 1, 23, 2, 0) op_5926 (v4740[22:0], v4741[17:0], v5926[22:0]); // 5.0
    wire [23:0] v5927; shift_adder #(24, 17, 1, 1, 24, 5, 0) op_5927 (v4742[23:0], v4743[16:0], v5927[23:0]); // 5.0
    wire [19:0] v5928; shift_adder #(19, 18, 1, 1, 20, 0, 0) op_5928 (v4744[18:0], v4623[17:0], v5928[19:0]); // 5.0
    wire [26:0] v5929; shift_adder #(16, 26, 1, 1, 27, -9, 0) op_5929 (v4745[15:0], v4746[25:0], v5929[26:0]); // 5.0
    wire [34:0] v5930; shift_adder #(35, 34, 1, 1, 35, 0, 0) op_5930 (v4747[34:0], v4748[33:0], v5930[34:0]); // 5.0
    wire [35:0] v5931; shift_adder #(27, 35, 1, 1, 36, -8, 0) op_5931 (v4749[26:0], v4750[34:0], v5931[35:0]); // 5.0
    wire [39:0] v5932; shift_adder #(39, 38, 1, 1, 40, 1, 0) op_5932 (v4751[38:0], v4752[37:0], v5932[39:0]); // 5.0
    wire [34:0] v5933; shift_adder #(35, 32, 1, 1, 35, 2, 0) op_5933 (v4753[34:0], v4754[31:0], v5933[34:0]); // 5.0
    wire [34:0] v5934; shift_adder #(34, 23, 1, 1, 35, 11, 0) op_5934 (v4690[33:0], v4755[22:0], v5934[34:0]); // 5.0
    wire [33:0] v5935; shift_adder #(29, 31, 1, 1, 34, -5, 0) op_5935 (v4756[28:0], v4663[30:0], v5935[33:0]); // 5.0
    wire [29:0] v5936; shift_adder #(25, 28, 1, 1, 30, -5, 0) op_5936 (v4757[24:0], v4758[27:0], v5936[29:0]); // 5.0
    wire [28:0] v5937; shift_adder #(29, 25, 1, 1, 29, 2, 0) op_5937 (v4759[28:0], v4760[24:0], v5937[28:0]); // 5.0
    wire [24:0] v5938; shift_adder #(23, 24, 1, 1, 25, -1, 0) op_5938 (v4761[22:0], v4762[23:0], v5938[24:0]); // 5.0
    wire [26:0] v5939; shift_adder #(8, 25, 1, 1, 27, 2, 0) op_5939 (v116[7:0], v4763[24:0], v5939[26:0]); // 5.0
    wire [25:0] v5940; shift_adder #(26, 21, 1, 1, 26, 4, 0) op_5940 (v4764[25:0], v4765[20:0], v5940[25:0]); // 5.0
    wire [24:0] v5941; shift_adder #(21, 25, 1, 1, 25, 0, 0) op_5941 (v4766[20:0], v4767[24:0], v5941[24:0]); // 5.0
    wire [24:0] v5942; shift_adder #(21, 24, 1, 1, 25, -2, 0) op_5942 (v4768[20:0], v4769[23:0], v5942[24:0]); // 5.0
    wire [28:0] v5943; shift_adder #(25, 29, 1, 1, 29, -3, 0) op_5943 (v4770[24:0], v4771[28:0], v5943[28:0]); // 5.0
    wire [22:0] v5944; shift_adder #(21, 21, 1, 1, 23, 2, 0) op_5944 (v4772[20:0], v4773[20:0], v5944[22:0]); // 5.0
    wire [32:0] v5945; shift_adder #(30, 33, 1, 1, 33, -1, 0) op_5945 (v4774[29:0], v4775[32:0], v5945[32:0]); // 5.0
    wire [34:0] v5946; shift_adder #(26, 33, 1, 1, 35, -8, 0) op_5946 (v4776[25:0], v4777[32:0], v5946[34:0]); // 5.0
    wire [33:0] v5947; shift_adder #(33, 25, 1, 1, 34, 9, 0) op_5947 (v4778[32:0], v4779[24:0], v5947[33:0]); // 5.0
    wire [38:0] v5948; shift_adder #(39, 15, 1, 1, 39, 2, 1) op_5948 (v4780[38:0], v4781[14:0], v5948[38:0]); // 5.0
    wire [19:0] v5949; shift_adder #(17, 18, 1, 1, 20, 2, 0) op_5949 (v4782[16:0], v4783[17:0], v5949[19:0]); // 5.0
    wire [30:0] v5950; shift_adder #(30, 23, 1, 1, 31, 8, 0) op_5950 (v4785[29:0], v4786[22:0], v5950[30:0]); // 5.0
    wire [18:0] v5951; shift_adder #(19, 16, 1, 1, 19, 0, 0) op_5951 (v4787[18:0], v4788[15:0], v5951[18:0]); // 5.0
    wire [21:0] v5952; shift_adder #(22, 18, 1, 1, 22, 2, 0) op_5952 (v4576[21:0], v4789[17:0], v5952[21:0]); // 5.0
    wire [27:0] v5953; shift_adder #(20, 26, 1, 1, 28, -7, 0) op_5953 (v4790[19:0], v4791[25:0], v5953[27:0]); // 5.0
    wire [24:0] v5954; shift_adder #(18, 24, 1, 1, 25, -6, 0) op_5954 (v4792[17:0], v4793[23:0], v5954[24:0]); // 5.0
    wire [17:0] v5955; shift_adder #(17, 15, 1, 1, 18, -1, 0) op_5955 (v4794[16:0], v4795[14:0], v5955[17:0]); // 5.0
    wire [24:0] v5956; shift_adder #(22, 23, 1, 1, 25, -2, 0) op_5956 (v4796[21:0], v4797[22:0], v5956[24:0]); // 5.0
    wire [26:0] v5957; shift_adder #(17, 26, 1, 1, 27, -8, 0) op_5957 (v4798[16:0], v4799[25:0], v5957[26:0]); // 5.0
    wire [28:0] v5958; shift_adder #(29, 25, 1, 1, 29, 2, 0) op_5958 (v4800[28:0], v4801[24:0], v5958[28:0]); // 5.0
    wire [29:0] v5959; shift_adder #(29, 29, 1, 1, 30, 0, 0) op_5959 (v4802[28:0], v4803[28:0], v5959[29:0]); // 5.0
    wire [26:0] v5960; shift_adder #(27, 25, 1, 1, 27, 0, 0) op_5960 (v4804[26:0], v4805[24:0], v5960[26:0]); // 5.0
    wire [28:0] v5961; shift_adder #(11, 22, 1, 1, 29, -18, 0) op_5961 (v153[10:0], v4806[21:0], v5961[28:0]); // 5.0
    wire [25:0] v5962; shift_adder #(8, 24, 1, 1, 26, 2, 0) op_5962 (v107[7:0], v4807[23:0], v5962[25:0]); // 5.0
    wire [28:0] v5963; shift_adder #(29, 20, 1, 1, 29, 7, 0) op_5963 (v4808[28:0], v4809[19:0], v5963[28:0]); // 5.0
    wire [22:0] v5964; shift_adder #(20, 20, 1, 1, 23, 2, 0) op_5964 (v4810[19:0], v4811[19:0], v5964[22:0]); // 5.0
    wire [27:0] v5965; shift_adder #(26, 26, 1, 1, 28, 1, 0) op_5965 (v4812[25:0], v4813[25:0], v5965[27:0]); // 5.0
    wire [28:0] v5966; shift_adder #(21, 28, 1, 1, 29, -7, 0) op_5966 (v4814[20:0], v4815[27:0], v5966[28:0]); // 5.0
    wire [25:0] v5967; shift_adder #(25, 19, 1, 1, 26, 4, 0) op_5967 (v4816[24:0], v4817[18:0], v5967[25:0]); // 5.0
    wire [25:0] v5968; shift_adder #(23, 24, 1, 1, 26, -2, 0) op_5968 (v4818[22:0], v4819[23:0], v5968[25:0]); // 5.0
    wire [23:0] v5969; shift_adder #(23, 20, 1, 1, 24, 1, 0) op_5969 (v4820[22:0], v4821[19:0], v5969[23:0]); // 5.0
    wire [25:0] v5970; shift_adder #(25, 19, 1, 1, 26, 4, 0) op_5970 (v4822[24:0], v4823[18:0], v5970[25:0]); // 5.0
    wire [22:0] v5971; shift_adder #(22, 19, 1, 1, 23, 1, 0) op_5971 (v4824[21:0], v4825[18:0], v5971[22:0]); // 5.0
    wire [21:0] v5972; shift_adder #(21, 20, 1, 1, 22, 1, 0) op_5972 (v4826[20:0], v4827[19:0], v5972[21:0]); // 5.0
    wire [24:0] v5973; shift_adder #(24, 21, 1, 1, 25, 3, 0) op_5973 (v4828[23:0], v4829[20:0], v5973[24:0]); // 5.0
    wire [22:0] v5974; shift_adder #(19, 23, 1, 1, 23, -1, 0) op_5974 (v4830[18:0], v4831[22:0], v5974[22:0]); // 5.0
    wire [25:0] v5975; shift_adder #(24, 25, 1, 1, 26, 0, 0) op_5975 (v4832[23:0], v4833[24:0], v5975[25:0]); // 5.0
    wire [29:0] v5976; shift_adder #(29, 26, 1, 1, 30, 3, 0) op_5976 (v4834[28:0], v4835[25:0], v5976[29:0]); // 5.0
    wire [23:0] v5977; shift_adder #(11, 24, 1, 1, 24, -8, 0) op_5977 (v287[10:0], v4836[23:0], v5977[23:0]); // 5.0
    wire [20:0] v5978; shift_adder #(16, 21, 1, 1, 21, -3, 0) op_5978 (v4837[15:0], v4838[20:0], v5978[20:0]); // 5.0
    wire [23:0] v5979; shift_adder #(20, 24, 1, 1, 24, -2, 0) op_5979 (v4840[19:0], v4841[23:0], v5979[23:0]); // 5.0
    wire [29:0] v5980; shift_adder #(27, 29, 1, 1, 30, -1, 0) op_5980 (v4842[26:0], v4843[28:0], v5980[29:0]); // 5.0
    wire [36:0] v5981; shift_adder #(18, 20, 1, 1, 37, 17, 1) op_5981 (v4844[17:0], v3188[19:0], v5981[36:0]); // 5.0
    wire [31:0] v5982; shift_adder #(31, 28, 1, 1, 32, 3, 0) op_5982 (v4845[30:0], v4846[27:0], v5982[31:0]); // 5.0
    wire [39:0] v5983; shift_adder #(39, 36, 1, 1, 40, 3, 0) op_5983 (v4847[38:0], v4848[35:0], v5983[39:0]); // 5.0
    wire [40:0] v5984; shift_adder #(25, 40, 1, 1, 41, -14, 0) op_5984 (v4849[24:0], v4850[39:0], v5984[40:0]); // 5.0
    wire [18:0] v5985; shift_adder #(18, 17, 1, 1, 19, 0, 0) op_5985 (v4851[17:0], v4852[16:0], v5985[18:0]); // 5.0
    wire [19:0] v5986; shift_adder #(18, 16, 1, 1, 20, 3, 0) op_5986 (v4853[17:0], v4854[15:0], v5986[19:0]); // 5.0
    wire [20:0] v5987; shift_adder #(20, 16, 1, 1, 21, 3, 0) op_5987 (v4855[19:0], v4856[15:0], v5987[20:0]); // 5.0
    wire [25:0] v5988; shift_adder #(20, 26, 1, 1, 26, -5, 0) op_5988 (v4857[19:0], v4858[25:0], v5988[25:0]); // 5.0
    wire [29:0] v5989; shift_adder #(26, 30, 1, 1, 30, -3, 0) op_5989 (v4859[25:0], v4860[29:0], v5989[29:0]); // 5.0
    wire [24:0] v5990; shift_adder #(19, 24, 1, 1, 25, -5, 0) op_5990 (v4861[18:0], v4862[23:0], v5990[24:0]); // 5.0
    wire [23:0] v5991; shift_adder #(21, 20, 1, 1, 24, 3, 0) op_5991 (v4863[20:0], v4864[19:0], v5991[23:0]); // 5.0
    wire [23:0] v5992; shift_adder #(22, 22, 1, 1, 24, -2, 0) op_5992 (v4865[21:0], v4866[21:0], v5992[23:0]); // 5.0
    wire [25:0] v5993; shift_adder #(23, 24, 1, 1, 26, -3, 0) op_5993 (v4867[22:0], v4868[23:0], v5993[25:0]); // 5.0
    wire [17:0] v5994; shift_adder #(11, 18, 1, 1, 18, -5, 0) op_5994 (v362[10:0], v4869[17:0], v5994[17:0]); // 5.0
    wire [34:0] v5995; shift_adder #(32, 26, 1, 1, 35, 9, 0) op_5995 (v4870[31:0], v4871[25:0], v5995[34:0]); // 5.0
    wire [26:0] v5996; shift_adder #(24, 26, 1, 1, 27, -2, 0) op_5996 (v4872[23:0], v4873[25:0], v5996[26:0]); // 5.0
    wire [19:0] v5997; shift_adder #(15, 19, 1, 1, 20, 1, 0) op_5997 (v4874[14:0], v4875[18:0], v5997[19:0]); // 5.0
    wire [38:0] v5998; shift_adder #(21, 38, 1, 1, 39, -15, 0) op_5998 (v4877[20:0], v4878[37:0], v5998[38:0]); // 5.0
    wire [31:0] v5999; shift_adder #(31, 26, 1, 1, 32, 5, 0) op_5999 (v4879[30:0], v4880[25:0], v5999[31:0]); // 5.0
    wire [34:0] v6000; shift_adder #(24, 34, 1, 1, 35, -11, 0) op_6000 (v4881[23:0], v4882[33:0], v6000[34:0]); // 5.0
    wire [32:0] v6001; shift_adder #(30, 32, 1, 1, 33, -3, 0) op_6001 (v4883[29:0], v4884[31:0], v6001[32:0]); // 5.0
    wire [29:0] v6002; shift_adder #(26, 29, 1, 1, 30, -3, 0) op_6002 (v4652[25:0], v4885[28:0], v6002[29:0]); // 5.0
    wire [29:0] v6003; shift_adder #(26, 28, 1, 1, 30, -3, 0) op_6003 (v4886[25:0], v4887[27:0], v6003[29:0]); // 5.0
    wire [32:0] v6004; shift_adder #(20, 31, 1, 1, 33, -13, 0) op_6004 (v4888[19:0], v4889[30:0], v6004[32:0]); // 5.0
    wire [25:0] v6005; shift_adder #(24, 24, 1, 1, 26, -2, 0) op_6005 (v4890[23:0], v4891[23:0], v6005[25:0]); // 5.0
    wire [22:0] v6006; shift_adder #(23, 22, 1, 1, 23, 0, 0) op_6006 (v4892[22:0], v4893[21:0], v6006[22:0]); // 5.0
    wire [23:0] v6007; shift_adder #(20, 20, 1, 1, 24, -4, 0) op_6007 (v4894[19:0], v4895[19:0], v6007[23:0]); // 5.0
    wire [22:0] v6008; shift_adder #(21, 22, 1, 1, 23, 1, 0) op_6008 (v4896[20:0], v4897[21:0], v6008[22:0]); // 5.0
    wire [20:0] v6009; shift_adder #(19, 16, 1, 1, 21, 4, 0) op_6009 (v4898[18:0], v4899[15:0], v6009[20:0]); // 5.0
    wire [22:0] v6010; shift_adder #(22, 18, 1, 1, 23, 4, 0) op_6010 (v4900[21:0], v4901[17:0], v6010[22:0]); // 5.0
    wire [25:0] v6011; shift_adder #(25, 20, 1, 1, 26, 6, 0) op_6011 (v4902[24:0], v4903[19:0], v6011[25:0]); // 5.0
    wire [35:0] v6012; shift_adder #(35, 19, 1, 1, 36, 15, 0) op_6012 (v4904[34:0], v4905[18:0], v6012[35:0]); // 5.0
    wire [30:0] v6013; shift_adder #(30, 19, 1, 1, 31, 11, 0) op_6013 (v4906[29:0], v4907[18:0], v6013[30:0]); // 5.0
    wire [34:0] v6014; shift_adder #(33, 23, 1, 1, 35, 12, 0) op_6014 (v4908[32:0], v4909[22:0], v6014[34:0]); // 5.0
    wire [28:0] v6015; shift_adder #(26, 29, 1, 1, 29, -1, 0) op_6015 (v4910[25:0], v4911[28:0], v6015[28:0]); // 5.0
    wire [30:0] v6016; shift_adder #(28, 22, 1, 1, 31, 9, 0) op_6016 (v4912[27:0], v4913[21:0], v6016[30:0]); // 5.0
    wire [36:0] v6017; shift_adder #(36, 33, 1, 1, 37, 3, 0) op_6017 (v4914[35:0], v4915[32:0], v6017[36:0]); // 5.0
    wire [39:0] v6018; shift_adder #(39, 34, 1, 1, 40, 5, 0) op_6018 (v4916[38:0], v4917[33:0], v6018[39:0]); // 5.0
    wire [37:0] v6019; shift_adder #(36, 37, 1, 1, 38, 0, 0) op_6019 (v4918[35:0], v4919[36:0], v6019[37:0]); // 5.0
    wire [23:0] v6020; shift_adder #(23, 20, 1, 1, 24, 1, 0) op_6020 (v4920[22:0], v4921[19:0], v6020[23:0]); // 5.0
    wire [19:0] v6021; shift_adder #(18, 18, 1, 1, 20, 2, 0) op_6021 (v4922[17:0], v4923[17:0], v6021[19:0]); // 5.0
    wire [33:0] v6022; shift_adder #(22, 33, 1, 1, 34, -11, 0) op_6022 (v4924[21:0], v4925[32:0], v6022[33:0]); // 5.0
    wire [31:0] v6023; shift_adder #(29, 31, 1, 1, 32, -3, 0) op_6023 (v4926[28:0], v4927[30:0], v6023[31:0]); // 5.0
    wire [31:0] v6024; shift_adder #(31, 29, 1, 1, 32, 3, 0) op_6024 (v4928[30:0], v4929[28:0], v6024[31:0]); // 5.0
    wire [26:0] v6025; shift_adder #(24, 25, 1, 1, 27, -2, 0) op_6025 (v4930[23:0], v4931[24:0], v6025[26:0]); // 5.0
    wire [26:0] v6026; shift_adder #(27, 25, 1, 1, 27, 1, 0) op_6026 (v4932[26:0], v4488[24:0], v6026[26:0]); // 5.0
    wire [30:0] v6027; shift_adder #(29, 28, 1, 1, 31, -2, 0) op_6027 (v4933[28:0], v4934[27:0], v6027[30:0]); // 5.0
    wire [23:0] v6028; shift_adder #(23, 20, 1, 1, 24, 4, 0) op_6028 (v4935[22:0], v4509[19:0], v6028[23:0]); // 5.0
    wire [22:0] v6029; shift_adder #(22, 20, 1, 1, 23, 2, 0) op_6029 (v4936[21:0], v4937[19:0], v6029[22:0]); // 5.0
    wire [28:0] v6030; shift_adder #(11, 25, 1, 1, 29, 4, 0) op_6030 (v145[10:0], v4938[24:0], v6030[28:0]); // 5.0
    wire [25:0] v6031; shift_adder #(20, 25, 1, 1, 26, -5, 0) op_6031 (v4939[19:0], v4940[24:0], v6031[25:0]); // 5.0
    wire [25:0] v6032; shift_adder #(24, 23, 1, 1, 26, 2, 0) op_6032 (v4671[23:0], v4941[22:0], v6032[25:0]); // 5.0
    wire [35:0] v6033; shift_adder #(32, 33, 1, 1, 36, -3, 0) op_6033 (v4942[31:0], v4943[32:0], v6033[35:0]); // 5.0
    wire [31:0] v6034; shift_adder #(32, 23, 1, 1, 32, 8, 0) op_6034 (v4944[31:0], v4945[22:0], v6034[31:0]); // 5.0
    wire [29:0] v6035; shift_adder #(24, 29, 1, 1, 30, -6, 0) op_6035 (v4819[23:0], v4946[28:0], v6035[29:0]); // 5.0
    wire [31:0] v6036; shift_adder #(26, 31, 1, 1, 32, -6, 0) op_6036 (v4947[25:0], v4948[30:0], v6036[31:0]); // 5.0
    wire [27:0] v6037; shift_adder #(28, 23, 1, 1, 28, 4, 0) op_6037 (v4949[27:0], v4950[22:0], v6037[27:0]); // 5.0
    wire [23:0] v6038; shift_adder #(23, 20, 1, 1, 24, 2, 0) op_6038 (v4951[22:0], v4952[19:0], v6038[23:0]); // 5.0
    wire [26:0] v6039; shift_adder #(26, 16, 1, 1, 27, 11, 0) op_6039 (v4953[25:0], v4954[15:0], v6039[26:0]); // 5.0
    wire [25:0] v6040; shift_adder #(23, 25, 1, 1, 26, -2, 0) op_6040 (v4955[22:0], v4956[24:0], v6040[25:0]); // 5.0
    wire [33:0] v6041; shift_adder #(24, 33, 1, 1, 34, -10, 0) op_6041 (v4957[23:0], v4958[32:0], v6041[33:0]); // 5.0
    wire [28:0] v6042; shift_adder #(10, 29, 1, 1, 29, -16, 1) op_6042 (v445[9:0], v4959[28:0], v6042[28:0]); // 5.0
    wire [30:0] v6043; shift_adder #(30, 26, 1, 1, 31, 3, 0) op_6043 (v4960[29:0], v4516[25:0], v6043[30:0]); // 5.0
    wire [19:0] v6044; shift_adder #(18, 19, 1, 1, 20, 1, 0) op_6044 (v4961[17:0], v4962[18:0], v6044[19:0]); // 5.0
    wire [31:0] v6045; shift_adder #(30, 24, 1, 1, 32, 8, 0) op_6045 (v4964[29:0], v4705[23:0], v6045[31:0]); // 5.0
    wire [34:0] v6046; shift_adder #(34, 34, 1, 1, 35, 0, 0) op_6046 (v4965[33:0], v4966[33:0], v6046[34:0]); // 5.0
    wire [38:0] v6047; shift_adder #(38, 25, 1, 1, 39, 13, 0) op_6047 (v4967[37:0], v4968[24:0], v6047[38:0]); // 5.0
    wire [35:0] v6048; shift_adder #(35, 19, 1, 1, 36, 16, 0) op_6048 (v4969[34:0], v4970[18:0], v6048[35:0]); // 5.0
    wire [39:0] v6049; shift_adder #(38, 17, 1, 1, 40, -2, 1) op_6049 (v4971[37:0], v4972[16:0], v6049[39:0]); // 5.0
    wire [20:0] v6050; shift_adder #(20, 17, 1, 1, 21, 2, 0) op_6050 (v4973[19:0], v4695[16:0], v6050[20:0]); // 5.0
    wire [22:0] v6051; shift_adder #(22, 22, 1, 1, 23, 0, 0) op_6051 (v4974[21:0], v4975[21:0], v6051[22:0]); // 5.0
    wire [25:0] v6052; shift_adder #(26, 17, 1, 1, 26, 5, 0) op_6052 (v4976[25:0], v4977[16:0], v6052[25:0]); // 5.0
    wire [19:0] v6053; shift_adder #(18, 19, 1, 1, 20, 1, 0) op_6053 (v4978[17:0], v4979[18:0], v6053[19:0]); // 5.0
    wire [25:0] v6054; shift_adder #(25, 22, 1, 1, 26, 4, 0) op_6054 (v4980[24:0], v4981[21:0], v6054[25:0]); // 5.0
    wire [29:0] v6055; shift_adder #(20, 29, 1, 1, 30, -9, 0) op_6055 (v4982[19:0], v4885[28:0], v6055[29:0]); // 5.0
    wire [30:0] v6056; shift_adder #(18, 30, 1, 1, 31, -11, 0) op_6056 (v4983[17:0], v4984[29:0], v6056[30:0]); // 5.0
    wire [30:0] v6057; shift_adder #(28, 30, 1, 1, 31, 1, 0) op_6057 (v4985[27:0], v4631[29:0], v6057[30:0]); // 5.0
    wire [27:0] v6058; shift_adder #(27, 19, 1, 1, 28, 9, 0) op_6058 (v4986[26:0], v4987[18:0], v6058[27:0]); // 5.0
    wire [28:0] v6059; shift_adder #(23, 28, 1, 1, 29, -4, 0) op_6059 (v4988[22:0], v4989[27:0], v6059[28:0]); // 5.0
    wire [36:0] v6060; shift_adder #(29, 36, 1, 1, 37, -6, 0) op_6060 (v4990[28:0], v4991[35:0], v6060[36:0]); // 5.0
    wire [20:0] v6061; shift_adder #(19, 17, 1, 1, 21, 3, 0) op_6061 (v4992[18:0], v4993[16:0], v6061[20:0]); // 5.0
    wire [30:0] v6062; shift_adder #(23, 30, 1, 1, 31, -6, 0) op_6062 (v4995[22:0], v4996[29:0], v6062[30:0]); // 5.0
    wire [38:0] v6063; shift_adder #(39, 14, 1, 1, 39, 3, 1) op_6063 (v4997[38:0], v4539[13:0], v6063[38:0]); // 5.0
    wire [25:0] v6064; shift_adder #(26, 17, 1, 1, 26, 7, 0) op_6064 (v4998[25:0], v4999[16:0], v6064[25:0]); // 5.0
    wire [22:0] v6065; shift_adder #(23, 19, 1, 1, 23, 2, 0) op_6065 (v5000[22:0], v5001[18:0], v6065[22:0]); // 5.0
    wire [20:0] v6066; shift_adder #(20, 18, 1, 1, 21, -1, 0) op_6066 (v5002[19:0], v5003[17:0], v6066[20:0]); // 5.0
    wire [19:0] v6067; shift_adder #(19, 17, 1, 1, 20, -1, 0) op_6067 (v5004[18:0], v5005[16:0], v6067[19:0]); // 5.0
    wire [27:0] v6068; shift_adder #(25, 26, 1, 1, 28, -2, 0) op_6068 (v5006[24:0], v5007[25:0], v6068[27:0]); // 5.0
    wire [26:0] v6069; shift_adder #(18, 26, 1, 1, 27, -8, 0) op_6069 (v5008[17:0], v5009[25:0], v6069[26:0]); // 5.0
    wire [25:0] v6070; shift_adder #(24, 24, 1, 1, 26, -1, 0) op_6070 (v5010[23:0], v5011[23:0], v6070[25:0]); // 5.0
    wire [31:0] v6071; shift_adder #(32, 28, 1, 1, 32, 2, 0) op_6071 (v4563[31:0], v5012[27:0], v6071[31:0]); // 5.0
    wire [31:0] v6072; shift_adder #(19, 29, 1, 1, 32, -13, 0) op_6072 (v5013[18:0], v4688[28:0], v6072[31:0]); // 5.0
    wire [29:0] v6073; shift_adder #(30, 25, 1, 1, 30, 3, 0) op_6073 (v5014[29:0], v5015[24:0], v6073[29:0]); // 5.0
    wire [26:0] v6074; shift_adder #(23, 26, 1, 1, 27, -2, 0) op_6074 (v4761[22:0], v5016[25:0], v6074[26:0]); // 5.0
    wire [26:0] v6075; shift_adder #(20, 26, 1, 1, 27, -5, 0) op_6075 (v5017[19:0], v5018[25:0], v6075[26:0]); // 5.0
    wire [21:0] v6076; shift_adder #(20, 18, 1, 1, 22, 4, 0) op_6076 (v5019[19:0], v5020[17:0], v6076[21:0]); // 5.0
    wire [26:0] v6077; shift_adder #(22, 26, 1, 1, 27, -3, 0) op_6077 (v5021[21:0], v5022[25:0], v6077[26:0]); // 5.0
    wire [22:0] v6078; shift_adder #(21, 20, 1, 1, 23, 3, 0) op_6078 (v5023[20:0], v5024[19:0], v6078[22:0]); // 5.0
    wire [22:0] v6079; shift_adder #(20, 19, 1, 1, 23, 4, 0) op_6079 (v5025[19:0], v5026[18:0], v6079[22:0]); // 5.0
    wire [29:0] v6080; shift_adder #(24, 29, 1, 1, 30, -5, 0) op_6080 (v5027[23:0], v5028[28:0], v6080[29:0]); // 5.0
    wire [27:0] v6081; shift_adder #(23, 28, 1, 1, 28, -3, 0) op_6081 (v4537[22:0], v5029[27:0], v6081[27:0]); // 5.0
    wire [33:0] v6082; shift_adder #(32, 27, 1, 1, 34, 6, 0) op_6082 (v4870[31:0], v5030[26:0], v6082[33:0]); // 5.0
    wire [28:0] v6083; shift_adder #(27, 20, 1, 1, 29, 8, 0) op_6083 (v5031[26:0], v5032[19:0], v6083[28:0]); // 5.0
    wire [40:0] v6084; shift_adder #(29, 41, 1, 1, 41, -11, 0) op_6084 (v4642[28:0], v5033[40:0], v6084[40:0]); // 5.0
    wire [33:0] v6085; shift_adder #(32, 15, 1, 1, 34, 18, 0) op_6085 (v5034[31:0], v5035[14:0], v6085[33:0]); // 5.0
    wire [27:0] v6086; shift_adder #(28, 19, 1, 1, 28, 7, 0) op_6086 (v5036[27:0], v5037[18:0], v6086[27:0]); // 5.0
    wire [21:0] v6087; shift_adder #(17, 19, 1, 1, 22, -4, 0) op_6087 (v5038[16:0], v5039[18:0], v6087[21:0]); // 5.0
    wire [20:0] v6088; shift_adder #(20, 21, 1, 1, 21, 0, 0) op_6088 (v5040[19:0], v5041[20:0], v6088[20:0]); // 5.0
    wire [37:0] v6089; shift_adder #(35, 38, 1, 1, 38, -2, 0) op_6089 (v5043[34:0], v5044[37:0], v6089[37:0]); // 5.0
    wire [18:0] v6090; shift_adder #(17, 17, 1, 1, 19, -1, 0) op_6090 (v5045[16:0], v5046[16:0], v6090[18:0]); // 5.0
    wire [34:0] v6091; shift_adder #(34, 15, 1, 1, 35, 18, 0) op_6091 (v5047[33:0], v5048[14:0], v6091[34:0]); // 5.0
    wire [24:0] v6092; shift_adder #(23, 24, 1, 1, 25, -1, 0) op_6092 (v5049[22:0], v5050[23:0], v6092[24:0]); // 5.0
    wire [33:0] v6093; shift_adder #(32, 33, 1, 1, 34, -2, 0) op_6093 (v5051[31:0], v4649[32:0], v6093[33:0]); // 5.0
    wire [29:0] v6094; shift_adder #(29, 27, 1, 1, 30, 1, 0) op_6094 (v5052[28:0], v5053[26:0], v6094[29:0]); // 5.0
    wire [29:0] v6095; shift_adder #(23, 29, 1, 1, 30, -6, 0) op_6095 (v5054[22:0], v5055[28:0], v6095[29:0]); // 5.0
    wire [30:0] v6096; shift_adder #(31, 20, 1, 1, 31, 9, 0) op_6096 (v5056[30:0], v5057[19:0], v6096[30:0]); // 5.0
    wire [26:0] v6097; shift_adder #(19, 25, 1, 1, 27, -7, 0) op_6097 (v5058[18:0], v5059[24:0], v6097[26:0]); // 5.0
    wire [22:0] v6098; shift_adder #(23, 16, 1, 1, 23, 4, 0) op_6098 (v5060[22:0], v4856[15:0], v6098[22:0]); // 5.0
    wire [25:0] v6099; shift_adder #(24, 17, 1, 1, 26, 9, 0) op_6099 (v5061[23:0], v5062[16:0], v6099[25:0]); // 5.0
    wire [22:0] v6100; shift_adder #(22, 19, 1, 1, 23, 3, 0) op_6100 (v5063[21:0], v5064[18:0], v6100[22:0]); // 5.0
    wire [23:0] v6101; shift_adder #(21, 22, 1, 1, 24, 2, 0) op_6101 (v5065[20:0], v4474[21:0], v6101[23:0]); // 5.0
    wire [27:0] v6102; shift_adder #(23, 18, 1, 1, 28, 10, 0) op_6102 (v5066[22:0], v5020[17:0], v6102[27:0]); // 5.0
    wire [32:0] v6103; shift_adder #(24, 33, 1, 1, 33, -6, 0) op_6103 (v5067[23:0], v5068[32:0], v6103[32:0]); // 5.0
    wire [26:0] v6104; shift_adder #(24, 23, 1, 1, 27, 3, 0) op_6104 (v5069[23:0], v5070[22:0], v6104[26:0]); // 5.0
    wire [33:0] v6105; shift_adder #(33, 25, 1, 1, 34, 8, 0) op_6105 (v5071[32:0], v5072[24:0], v6105[33:0]); // 5.0
    wire [39:0] v6106; shift_adder #(25, 39, 1, 1, 40, -14, 0) op_6106 (v5073[24:0], v5074[38:0], v6106[39:0]); // 5.0
    wire [40:0] v6107; shift_adder #(41, 19, 1, 1, 41, 0, 1) op_6107 (v5075[40:0], v5076[18:0], v6107[40:0]); // 5.0
    wire [25:0] v6108; shift_adder #(26, 17, 1, 1, 26, 6, 0) op_6108 (v5077[25:0], v5078[16:0], v6108[25:0]); // 5.0
    wire [21:0] v6109; shift_adder #(18, 20, 1, 1, 22, -4, 0) op_6109 (v5079[17:0], v5080[19:0], v6109[21:0]); // 5.0
    wire [18:0] v6110; shift_adder #(16, 18, 1, 1, 19, -1, 0) op_6110 (v5081[15:0], v5082[17:0], v6110[18:0]); // 5.0
    wire [36:0] v6111; shift_adder #(36, 22, 1, 1, 37, 14, 0) op_6111 (v5084[35:0], v5085[21:0], v6111[36:0]); // 5.0
    wire [18:0] v6112; shift_adder #(19, 16, 1, 1, 19, 0, 0) op_6112 (v5086[18:0], v5087[15:0], v6112[18:0]); // 5.0
    wire [33:0] v6113; shift_adder #(32, 34, 1, 1, 34, -1, 0) op_6113 (v5088[31:0], v5089[33:0], v6113[33:0]); // 5.0
    wire [33:0] v6114; shift_adder #(34, 28, 1, 1, 34, 5, 0) op_6114 (v5090[33:0], v5091[27:0], v6114[33:0]); // 5.0
    wire [30:0] v6115; shift_adder #(29, 30, 1, 1, 31, 0, 0) op_6115 (v5092[28:0], v5093[29:0], v6115[30:0]); // 5.0
    wire [32:0] v6116; shift_adder #(33, 31, 1, 1, 33, 0, 0) op_6116 (v5094[32:0], v4646[30:0], v6116[32:0]); // 5.0
    wire [26:0] v6117; shift_adder #(25, 26, 1, 1, 27, -2, 0) op_6117 (v5095[24:0], v5096[25:0], v6117[26:0]); // 5.0
    wire [30:0] v6118; shift_adder #(8, 26, 1, 1, 31, 5, 1) op_6118 (v79[7:0], v5097[25:0], v6118[30:0]); // 5.0
    wire [23:0] v6119; shift_adder #(23, 21, 1, 1, 24, 1, 0) op_6119 (v5098[22:0], v5099[20:0], v6119[23:0]); // 5.0
    wire [28:0] v6120; shift_adder #(29, 22, 1, 1, 29, 5, 0) op_6120 (v5100[28:0], v5101[21:0], v6120[28:0]); // 5.0
    wire [30:0] v6121; shift_adder #(26, 30, 1, 1, 31, -4, 0) op_6121 (v5102[25:0], v5103[29:0], v6121[30:0]); // 5.0
    wire [29:0] v6122; shift_adder #(30, 20, 1, 1, 30, 9, 0) op_6122 (v5104[29:0], v4903[19:0], v6122[29:0]); // 5.0
    wire [26:0] v6123; shift_adder #(26, 20, 1, 1, 27, 6, 0) op_6123 (v5105[25:0], v5106[19:0], v6123[26:0]); // 5.0
    wire [26:0] v6124; shift_adder #(26, 16, 1, 1, 27, 11, 0) op_6124 (v5107[25:0], v5108[15:0], v6124[26:0]); // 5.0
    wire [22:0] v6125; shift_adder #(21, 23, 1, 1, 23, -1, 0) op_6125 (v5109[20:0], v5110[22:0], v6125[22:0]); // 5.0
    wire [26:0] v6126; shift_adder #(25, 27, 1, 1, 27, 0, 0) op_6126 (v5111[24:0], v5112[26:0], v6126[26:0]); // 5.0
    wire [26:0] v6127; shift_adder #(15, 26, 1, 1, 27, -12, 0) op_6127 (v5113[14:0], v5114[25:0], v6127[26:0]); // 5.0
    wire [20:0] v6128; shift_adder #(17, 21, 1, 1, 21, -1, 0) op_6128 (v5115[16:0], v5116[20:0], v6128[20:0]); // 5.0
    wire [36:0] v6129; shift_adder #(17, 31, 1, 1, 37, 6, 1) op_6129 (v5118[16:0], v3605[30:0], v6129[36:0]); // 5.0
    wire [34:0] v6130; shift_adder #(34, 29, 1, 1, 35, 5, 0) op_6130 (v5119[33:0], v5120[28:0], v6130[34:0]); // 5.0
    wire [37:0] v6131; shift_adder #(24, 37, 1, 1, 38, -13, 0) op_6131 (v5121[23:0], v5122[36:0], v6131[37:0]); // 5.0
    wire [41:0] v6132; shift_adder #(41, 38, 1, 1, 42, 3, 0) op_6132 (v5123[40:0], v5124[37:0], v6132[41:0]); // 5.0
    wire [20:0] v6133; shift_adder #(20, 16, 1, 1, 21, 3, 0) op_6133 (v5125[19:0], v4745[15:0], v6133[20:0]); // 5.0
    wire [18:0] v6134; shift_adder #(17, 16, 1, 1, 19, -1, 0) op_6134 (v5126[16:0], v5127[15:0], v6134[18:0]); // 5.0
    wire [25:0] v6135; shift_adder #(25, 23, 1, 1, 26, 2, 0) op_6135 (v5128[24:0], v5129[22:0], v6135[25:0]); // 5.0
    wire [29:0] v6136; shift_adder #(29, 25, 1, 1, 30, 3, 0) op_6136 (v5130[28:0], v5131[24:0], v6136[29:0]); // 5.0
    wire [29:0] v6137; shift_adder #(25, 28, 1, 1, 30, -4, 0) op_6137 (v5132[24:0], v5133[27:0], v6137[29:0]); // 5.0
    wire [26:0] v6138; shift_adder #(26, 19, 1, 1, 27, 6, 0) op_6138 (v5134[25:0], v5135[18:0], v6138[26:0]); // 5.0
    wire [26:0] v6139; shift_adder #(22, 26, 1, 1, 27, -4, 0) op_6139 (v4491[21:0], v5136[25:0], v6139[26:0]); // 5.0
    wire [26:0] v6140; shift_adder #(25, 25, 1, 1, 27, -1, 0) op_6140 (v5137[24:0], v5138[24:0], v6140[26:0]); // 5.0
    wire [24:0] v6141; shift_adder #(23, 23, 1, 1, 25, -1, 0) op_6141 (v5139[22:0], v5140[22:0], v6141[24:0]); // 5.0
    wire [23:0] v6142; shift_adder #(17, 22, 1, 1, 24, -6, 0) op_6142 (v5141[16:0], v5142[21:0], v6142[23:0]); // 5.0
    wire [21:0] v6143; shift_adder #(11, 19, 1, 1, 22, 3, 1) op_6143 (v659[10:0], v5143[18:0], v6143[21:0]); // 5.0
    wire [22:0] v6144; shift_adder #(22, 22, 1, 1, 23, 0, 0) op_6144 (v5144[21:0], v5145[21:0], v6144[22:0]); // 5.0
    wire [25:0] v6145; shift_adder #(23, 22, 1, 1, 26, 3, 0) op_6145 (v5146[22:0], v5147[21:0], v6145[25:0]); // 5.0
    wire [31:0] v6146; shift_adder #(30, 26, 1, 1, 32, 5, 0) op_6146 (v5148[29:0], v5149[25:0], v6146[31:0]); // 5.0
    wire [21:0] v6147; shift_adder #(22, 19, 1, 1, 22, 2, 0) op_6147 (v5150[21:0], v5151[18:0], v6147[21:0]); // 5.0
    wire [35:0] v6148; shift_adder #(29, 35, 1, 1, 36, -6, 0) op_6148 (v5152[28:0], v5153[34:0], v6148[35:0]); // 5.0
    wire [26:0] v6149; shift_adder #(19, 25, 1, 1, 27, -8, 0) op_6149 (v5154[18:0], v5155[24:0], v6149[26:0]); // 5.0
    wire [31:0] v6150; shift_adder #(16, 31, 1, 1, 32, -14, 0) op_6150 (v5156[15:0], v5157[30:0], v6150[31:0]); // 5.0
    wire [35:0] v6151; shift_adder #(34, 20, 1, 1, 36, 15, 0) op_6151 (v5158[33:0], v5159[19:0], v6151[35:0]); // 5.0
    wire [18:0] v6152; shift_adder #(15, 17, 1, 1, 19, -3, 0) op_6152 (v5160[14:0], v5161[16:0], v6152[18:0]); // 5.0
    wire [19:0] v6153; shift_adder #(20, 18, 1, 1, 20, 0, 0) op_6153 (v5162[19:0], v5163[17:0], v6153[19:0]); // 5.0
    wire [19:0] v6154; shift_adder #(20, 17, 1, 1, 20, 0, 0) op_6154 (v5164[19:0], v5165[16:0], v6154[19:0]); // 5.0
    wire [26:0] v6155; shift_adder #(18, 27, 1, 1, 27, -8, 0) op_6155 (v5166[17:0], v5167[26:0], v6155[26:0]); // 5.0
    wire [28:0] v6156; shift_adder #(26, 27, 1, 1, 29, -2, 0) op_6156 (v5168[25:0], v5169[26:0], v6156[28:0]); // 5.0
    wire [22:0] v6157; shift_adder #(20, 21, 1, 1, 23, -2, 0) op_6157 (v5170[19:0], v5171[20:0], v6157[22:0]); // 5.0
    wire [28:0] v6158; shift_adder #(25, 26, 1, 1, 29, -3, 0) op_6158 (v5172[24:0], v5173[25:0], v6158[28:0]); // 5.0
    wire [30:0] v6159; shift_adder #(26, 31, 1, 1, 31, -1, 0) op_6159 (v5174[25:0], v5175[30:0], v6159[30:0]); // 5.0
    wire [32:0] v6160; shift_adder #(31, 22, 1, 1, 33, 10, 0) op_6160 (v5176[30:0], v5177[21:0], v6160[32:0]); // 5.0
    wire [32:0] v6161; shift_adder #(27, 33, 1, 1, 33, -4, 0) op_6161 (v5178[26:0], v5179[32:0], v6161[32:0]); // 5.0
    wire [20:0] v6162; shift_adder #(18, 19, 1, 1, 21, 2, 0) op_6162 (v5180[17:0], v5181[18:0], v6162[20:0]); // 5.0
    wire [35:0] v6163; shift_adder #(34, 25, 1, 1, 36, 10, 0) op_6163 (v5183[33:0], v4602[24:0], v6163[35:0]); // 5.0
    wire [33:0] v6164; shift_adder #(15, 24, 1, 1, 34, 10, 1) op_6164 (v5184[14:0], v3379[23:0], v6164[33:0]); // 5.0
    wire [25:0] v6165; shift_adder #(18, 26, 1, 1, 26, -7, 0) op_6165 (v5185[17:0], v5186[25:0], v6165[25:0]); // 5.0
    wire [25:0] v6166; shift_adder #(24, 23, 1, 1, 26, 2, 0) op_6166 (v5187[23:0], v5188[22:0], v6166[25:0]); // 5.0
    wire [26:0] v6167; shift_adder #(25, 16, 1, 1, 27, 10, 0) op_6167 (v4464[24:0], v5189[15:0], v6167[26:0]); // 5.0
    wire [28:0] v6168; shift_adder #(27, 28, 1, 1, 29, 0, 0) op_6168 (v5190[26:0], v5191[27:0], v6168[28:0]); // 5.0
    wire [27:0] v6169; shift_adder #(19, 27, 1, 1, 28, -9, 0) op_6169 (v5192[18:0], v5193[26:0], v6169[27:0]); // 5.0
    wire [23:0] v6170; shift_adder #(23, 22, 1, 1, 24, 1, 0) op_6170 (v5194[22:0], v5195[21:0], v6170[23:0]); // 5.0
    wire [34:0] v6171; shift_adder #(34, 14, 1, 1, 35, 19, 0) op_6171 (v5196[33:0], v5197[13:0], v6171[34:0]); // 5.0
    wire [27:0] v6172; shift_adder #(25, 27, 1, 1, 28, -2, 0) op_6172 (v5198[24:0], v5199[26:0], v6172[27:0]); // 5.0
    wire [32:0] v6173; shift_adder #(12, 27, 1, 1, 33, 6, 1) op_6173 (v2033[11:0], v5200[26:0], v6173[32:0]); // 5.0
    wire [19:0] v6174; shift_adder #(19, 16, 1, 1, 20, 3, 0) op_6174 (v5201[18:0], v5202[15:0], v6174[19:0]); // 5.0
    wire [20:0] v6175; shift_adder #(19, 21, 1, 1, 21, 0, 0) op_6175 (v5203[18:0], v5204[20:0], v6175[20:0]); // 5.0
    wire [36:0] v6176; shift_adder #(23, 35, 1, 1, 37, -13, 0) op_6176 (v5205[22:0], v5206[34:0], v6176[36:0]); // 5.0
    wire [28:0] v6177; shift_adder #(28, 25, 1, 1, 29, 3, 0) op_6177 (v5207[27:0], v5208[24:0], v6177[28:0]); // 5.0
    wire [19:0] v6178; shift_adder #(18, 18, 1, 1, 20, -1, 0) op_6178 (v5209[17:0], v5210[17:0], v6178[19:0]); // 5.0
    wire [25:0] v6179; shift_adder #(24, 20, 1, 1, 26, 5, 0) op_6179 (v5211[23:0], v5162[19:0], v6179[25:0]); // 5.0
    wire [25:0] v6180; shift_adder #(26, 21, 1, 1, 26, 4, 0) op_6180 (v5212[25:0], v5213[20:0], v6180[25:0]); // 5.0
    wire [25:0] v6181; shift_adder #(20, 26, 1, 1, 26, -3, 0) op_6181 (v5214[19:0], v5215[25:0], v6181[25:0]); // 5.0
    wire [38:0] v6182; shift_adder #(38, 24, 1, 1, 39, 13, 0) op_6182 (v5216[37:0], v5217[23:0], v6182[38:0]); // 5.0
    wire [25:0] v6183; shift_adder #(15, 25, 1, 1, 26, -9, 0) op_6183 (v4719[14:0], v5218[24:0], v6183[25:0]); // 5.0
    wire [35:0] v6184; shift_adder #(34, 31, 1, 1, 36, 4, 0) op_6184 (v5219[33:0], v5220[30:0], v6184[35:0]); // 5.0
    wire [38:0] v6185; shift_adder #(38, 17, 1, 1, 39, -1, 1) op_6185 (v5221[37:0], v5222[16:0], v6185[38:0]); // 5.0
    wire [18:0] v6186; shift_adder #(17, 16, 1, 1, 19, -1, 0) op_6186 (v5223[16:0], v5224[15:0], v6186[18:0]); // 5.0
    wire [21:0] v6187; shift_adder #(21, 20, 1, 1, 22, 1, 0) op_6187 (v5225[20:0], v5226[19:0], v6187[21:0]); // 5.0
    wire [21:0] v6188; shift_adder #(21, 21, 1, 1, 22, -1, 0) op_6188 (v5227[20:0], v5228[20:0], v6188[21:0]); // 5.0
    wire [23:0] v6189; shift_adder #(19, 23, 1, 1, 24, -3, 0) op_6189 (v5229[18:0], v5230[22:0], v6189[23:0]); // 5.0
    wire [24:0] v6190; shift_adder #(23, 24, 1, 1, 25, 0, 0) op_6190 (v5231[22:0], v5232[23:0], v6190[24:0]); // 5.0
    wire [26:0] v6191; shift_adder #(22, 26, 1, 1, 27, -3, 0) op_6191 (v5233[21:0], v5234[25:0], v6191[26:0]); // 5.0
    wire [26:0] v6192; shift_adder #(26, 26, 1, 1, 27, 0, 0) op_6192 (v5235[25:0], v4506[25:0], v6192[26:0]); // 5.0
    wire [30:0] v6193; shift_adder #(25, 30, 1, 1, 31, -4, 0) op_6193 (v5236[24:0], v5237[29:0], v6193[30:0]); // 5.0
    wire [28:0] v6194; shift_adder #(28, 19, 1, 1, 29, 10, 0) op_6194 (v5238[27:0], v4650[18:0], v6194[28:0]); // 5.0
    wire [30:0] v6195; shift_adder #(29, 26, 1, 1, 31, 4, 0) op_6195 (v5239[28:0], v5240[25:0], v6195[30:0]); // 5.0
    wire [18:0] v6196; shift_adder #(18, 16, 1, 1, 19, 2, 0) op_6196 (v5241[17:0], v5242[15:0], v6196[18:0]); // 5.0
    wire [23:0] v6197; shift_adder #(23, 21, 1, 1, 24, 0, 0) op_6197 (v5244[22:0], v5245[20:0], v6197[23:0]); // 5.0
    wire [20:0] v6198; shift_adder #(21, 15, 1, 1, 21, 1, 0) op_6198 (v5246[20:0], v5247[14:0], v6198[20:0]); // 5.0
    wire [32:0] v6199; shift_adder #(32, 30, 1, 1, 33, 2, 0) op_6199 (v5248[31:0], v5249[29:0], v6199[32:0]); // 5.0
    wire [35:0] v6200; shift_adder #(36, 14, 1, 1, 36, 2, 1) op_6200 (v5250[35:0], v5197[13:0], v6200[35:0]); // 5.0
    wire [36:0] v6201; shift_adder #(36, 25, 1, 1, 37, 11, 0) op_6201 (v5251[35:0], v5252[24:0], v6201[36:0]); // 5.0
    wire [38:0] v6202; shift_adder #(38, 34, 1, 1, 39, 3, 0) op_6202 (v5253[37:0], v5254[33:0], v6202[38:0]); // 5.0
    wire [29:0] v6203; shift_adder #(24, 30, 1, 1, 30, -5, 0) op_6203 (v5255[23:0], v5256[29:0], v6203[29:0]); // 5.0
    wire [27:0] v6204; shift_adder #(27, 17, 1, 1, 28, 10, 0) op_6204 (v5257[26:0], v5258[16:0], v6204[27:0]); // 5.0
    wire [27:0] v6205; shift_adder #(28, 17, 1, 1, 28, 8, 0) op_6205 (v5259[27:0], v5260[16:0], v6205[27:0]); // 5.0
    wire [29:0] v6206; shift_adder #(26, 30, 1, 1, 30, -3, 0) op_6206 (v5261[25:0], v5262[29:0], v6206[29:0]); // 5.0
    wire [30:0] v6207; shift_adder #(27, 29, 1, 1, 31, -3, 0) op_6207 (v5263[26:0], v5264[28:0], v6207[30:0]); // 5.0
    wire [25:0] v6208; shift_adder #(25, 18, 1, 1, 26, 7, 0) op_6208 (v5265[24:0], v5266[17:0], v6208[25:0]); // 5.0
    wire [24:0] v6209; shift_adder #(11, 23, 1, 1, 25, -14, 1) op_6209 (v188[10:0], v5267[22:0], v6209[24:0]); // 5.0
    wire [26:0] v6210; shift_adder #(18, 25, 1, 1, 27, -9, 0) op_6210 (v4789[17:0], v5268[24:0], v6210[26:0]); // 5.0
    wire [25:0] v6211; shift_adder #(23, 20, 1, 1, 26, 6, 0) op_6211 (v5269[22:0], v4526[19:0], v6211[25:0]); // 5.0
    wire [20:0] v6212; shift_adder #(18, 20, 1, 1, 21, -2, 0) op_6212 (v5270[17:0], v5271[19:0], v6212[20:0]); // 5.0
    wire [24:0] v6213; shift_adder #(22, 25, 1, 1, 25, -1, 0) op_6213 (v5272[21:0], v5273[24:0], v6213[24:0]); // 5.0
    wire [25:0] v6214; shift_adder #(21, 25, 1, 1, 26, -3, 0) op_6214 (v5274[20:0], v5275[24:0], v6214[25:0]); // 5.0
    wire [27:0] v6215; shift_adder #(26, 25, 1, 1, 28, 3, 0) op_6215 (v5276[25:0], v5277[24:0], v6215[27:0]); // 5.0
    wire [27:0] v6216; shift_adder #(26, 27, 1, 1, 28, -2, 0) op_6216 (v5278[25:0], v5279[26:0], v6216[27:0]); // 5.0
    wire [32:0] v6217; shift_adder #(26, 32, 1, 1, 33, -6, 0) op_6217 (v5280[25:0], v5281[31:0], v6217[32:0]); // 5.0
    wire [30:0] v6218; shift_adder #(24, 31, 1, 1, 31, -4, 0) op_6218 (v5282[23:0], v5283[30:0], v6218[30:0]); // 5.0
    wire [36:0] v6219; shift_adder #(37, 16, 1, 1, 37, 0, 1) op_6219 (v5284[36:0], v5285[15:0], v6219[36:0]); // 5.0
    wire [39:0] v6220; shift_adder #(39, 39, 1, 1, 40, 0, 0) op_6220 (v5286[38:0], v5287[38:0], v6220[39:0]); // 5.0
    wire [24:0] v6221; shift_adder #(24, 23, 1, 1, 25, -1, 0) op_6221 (v5288[23:0], v5289[22:0], v6221[24:0]); // 5.0
    wire [18:0] v6222; shift_adder #(17, 17, 1, 1, 19, -1, 0) op_6222 (v5290[16:0], v5291[16:0], v6222[18:0]); // 5.0
    wire [20:0] v6223; shift_adder #(19, 19, 1, 1, 21, 2, 0) op_6223 (v5292[18:0], v5293[18:0], v6223[20:0]); // 5.0
    wire [33:0] v6224; shift_adder #(33, 23, 1, 1, 34, 10, 0) op_6224 (v5295[32:0], v5296[22:0], v6224[33:0]); // 5.0
    wire [27:0] v6225; shift_adder #(27, 20, 1, 1, 28, 7, 0) op_6225 (v5297[26:0], v5298[19:0], v6225[27:0]); // 5.0
    wire [28:0] v6226; shift_adder #(28, 24, 1, 1, 29, 4, 0) op_6226 (v5299[27:0], v5300[23:0], v6226[28:0]); // 5.0
    wire [32:0] v6227; shift_adder #(29, 31, 1, 1, 33, -3, 0) op_6227 (v5301[28:0], v4845[30:0], v6227[32:0]); // 5.0
    wire [34:0] v6228; shift_adder #(32, 33, 1, 1, 35, -3, 0) op_6228 (v5302[31:0], v5303[32:0], v6228[34:0]); // 5.0
    wire [34:0] v6229; shift_adder #(25, 33, 1, 1, 35, -9, 0) op_6229 (v5304[24:0], v5305[32:0], v6229[34:0]); // 5.0
    wire [24:0] v6230; shift_adder #(18, 23, 1, 1, 25, -7, 0) op_6230 (v5306[17:0], v5307[22:0], v6230[24:0]); // 5.0
    wire [27:0] v6231; shift_adder #(27, 26, 1, 1, 28, -1, 0) op_6231 (v5308[26:0], v5309[25:0], v6231[27:0]); // 5.0
    wire [30:0] v6232; shift_adder #(30, 22, 1, 1, 31, 8, 0) op_6232 (v5310[29:0], v5311[21:0], v6232[30:0]); // 5.0
    wire [24:0] v6233; shift_adder #(23, 18, 1, 1, 25, 6, 0) op_6233 (v5312[22:0], v5313[17:0], v6233[24:0]); // 5.0
    wire [27:0] v6234; shift_adder #(21, 27, 1, 1, 28, -5, 0) op_6234 (v5314[20:0], v5315[26:0], v6234[27:0]); // 5.0
    wire [36:0] v6235; shift_adder #(28, 35, 1, 1, 37, -8, 0) op_6235 (v5316[27:0], v5317[34:0], v6235[36:0]); // 5.0
    wire [19:0] v6236; shift_adder #(18, 18, 1, 1, 20, 2, 0) op_6236 (v5318[17:0], v5319[17:0], v6236[19:0]); // 5.0
    wire [26:0] v6237; shift_adder #(25, 19, 1, 1, 27, 7, 0) op_6237 (v5320[24:0], v5321[18:0], v6237[26:0]); // 5.0
    wire [36:0] v6238; shift_adder #(36, 23, 1, 1, 37, 13, 0) op_6238 (v5322[35:0], v5323[22:0], v6238[36:0]); // 5.0
    wire [33:0] v6239; shift_adder #(15, 17, 1, 1, 34, 17, 1) op_6239 (v4710[14:0], v3889[16:0], v6239[33:0]); // 5.0
    wire [32:0] v6240; shift_adder #(32, 31, 1, 1, 33, 1, 0) op_6240 (v5324[31:0], v4626[30:0], v6240[32:0]); // 5.0
    wire [28:0] v6241; shift_adder #(28, 21, 1, 1, 29, 7, 0) op_6241 (v5325[27:0], v5326[20:0], v6241[28:0]); // 5.0
    wire [39:0] v6242; shift_adder #(30, 39, 1, 1, 40, -8, 0) op_6242 (v5327[29:0], v5328[38:0], v6242[39:0]); // 5.0
    wire [38:0] v6243; shift_adder #(37, 37, 1, 1, 39, 1, 0) op_6243 (v5329[36:0], v5330[36:0], v6243[38:0]); // 5.0
    wire [21:0] v6244; shift_adder #(21, 19, 1, 1, 22, 0, 0) op_6244 (v5331[20:0], v5332[18:0], v6244[21:0]); // 5.0
    wire [20:0] v6245; shift_adder #(16, 19, 1, 1, 21, -5, 0) op_6245 (v5333[15:0], v5334[18:0], v6245[20:0]); // 5.0
    wire [35:0] v6246; shift_adder #(21, 34, 1, 1, 36, -14, 0) op_6246 (v5335[20:0], v5336[33:0], v6246[35:0]); // 5.0
    wire [32:0] v6247; shift_adder #(27, 32, 1, 1, 33, -5, 0) op_6247 (v5337[26:0], v5338[31:0], v6247[32:0]); // 5.0
    wire [28:0] v6248; shift_adder #(22, 26, 1, 1, 29, -7, 0) op_6248 (v5339[21:0], v5340[25:0], v6248[28:0]); // 5.0
    wire [22:0] v6249; shift_adder #(18, 23, 1, 1, 23, -3, 0) op_6249 (v5341[17:0], v5342[22:0], v6249[22:0]); // 5.0
    wire [21:0] v6250; shift_adder #(19, 18, 1, 1, 22, -2, 0) op_6250 (v5343[18:0], v5344[17:0], v6250[21:0]); // 5.0
    wire [22:0] v6251; shift_adder #(21, 22, 1, 1, 23, -1, 0) op_6251 (v5225[20:0], v5345[21:0], v6251[22:0]); // 5.0
    wire [23:0] v6252; shift_adder #(22, 23, 1, 1, 24, -1, 0) op_6252 (v5346[21:0], v5342[22:0], v6252[23:0]); // 5.0
    wire [21:0] v6253; shift_adder #(17, 21, 1, 1, 22, -4, 0) op_6253 (v5347[16:0], v5348[20:0], v6253[21:0]); // 5.0
    wire [20:0] v6254; shift_adder #(19, 20, 1, 1, 21, -1, 0) op_6254 (v5349[18:0], v5350[19:0], v6254[20:0]); // 5.0
    wire [29:0] v6255; shift_adder #(25, 30, 1, 1, 30, -2, 0) op_6255 (v5351[24:0], v5352[29:0], v6255[29:0]); // 5.0
    wire [28:0] v6256; shift_adder #(27, 23, 1, 1, 29, 6, 0) op_6256 (v5257[26:0], v5353[22:0], v6256[28:0]); // 5.0
    wire [22:0] v6257; shift_adder #(21, 18, 1, 1, 23, 5, 0) op_6257 (v5354[20:0], v5355[17:0], v6257[22:0]); // 5.0
    wire [26:0] v6258; shift_adder #(24, 26, 1, 1, 27, 1, 0) op_6258 (v4645[23:0], v5356[25:0], v6258[26:0]); // 5.0
    wire [31:0] v6259; shift_adder #(22, 31, 1, 1, 32, -8, 0) op_6259 (v5357[21:0], v5358[30:0], v6259[31:0]); // 5.0
    wire [18:0] v6260; shift_adder #(15, 19, 1, 1, 19, -1, 0) op_6260 (v5359[14:0], v5360[18:0], v6260[18:0]); // 5.0
    wire [39:0] v6261; shift_adder #(40, 23, 1, 1, 40, 16, 0) op_6261 (v5362[39:0], v5363[22:0], v6261[39:0]); // 5.0
    wire [36:0] v6262; shift_adder #(37, 14, 1, 1, 37, 1, 1) op_6262 (v5364[36:0], v5365[13:0], v6262[36:0]); // 5.0
    wire [26:0] v6263; shift_adder #(26, 17, 1, 1, 27, 8, 0) op_6263 (v5366[25:0], v5367[16:0], v6263[26:0]); // 5.0
    wire [21:0] v6264; shift_adder #(8, 20, 1, 1, 22, 2, 1) op_6264 (v66[7:0], v5368[19:0], v6264[21:0]); // 5.0
    wire [22:0] v6265; shift_adder #(21, 22, 1, 1, 23, 1, 0) op_6265 (v5369[20:0], v4726[21:0], v6265[22:0]); // 5.0
    wire [19:0] v6266; shift_adder #(18, 18, 1, 1, 20, -1, 0) op_6266 (v5370[17:0], v5371[17:0], v6266[19:0]); // 5.0
    wire [30:0] v6267; shift_adder #(22, 29, 1, 1, 31, -9, 0) op_6267 (v5372[21:0], v5373[28:0], v6267[30:0]); // 5.0
    wire [24:0] v6268; shift_adder #(16, 23, 1, 1, 25, -8, 0) op_6268 (v5374[15:0], v5375[22:0], v6268[24:0]); // 5.0
    wire [18:0] v6269; shift_adder #(18, 17, 1, 1, 19, 1, 0) op_6269 (v5376[17:0], v5377[16:0], v6269[18:0]); // 5.0
    wire [29:0] v6270; shift_adder #(29, 24, 1, 1, 30, 3, 0) op_6270 (v5378[28:0], v5379[23:0], v6270[29:0]); // 5.0
    wire [29:0] v6271; shift_adder #(30, 25, 1, 1, 30, 1, 0) op_6271 (v5380[29:0], v5381[24:0], v6271[29:0]); // 5.0
    wire [28:0] v6272; shift_adder #(28, 22, 1, 1, 29, 5, 0) op_6272 (v5382[27:0], v4732[21:0], v6272[28:0]); // 5.0
    wire [24:0] v6273; shift_adder #(17, 23, 1, 1, 25, -7, 0) op_6273 (v5383[16:0], v5384[22:0], v6273[24:0]); // 5.0
    wire [22:0] v6274; shift_adder #(19, 21, 1, 1, 23, 2, 0) op_6274 (v5385[18:0], v5386[20:0], v6274[22:0]); // 5.0
    wire [26:0] v6275; shift_adder #(26, 21, 1, 1, 27, 4, 0) op_6275 (v5387[25:0], v5388[20:0], v6275[26:0]); // 5.0
    wire [24:0] v6276; shift_adder #(17, 25, 1, 1, 25, -7, 0) op_6276 (v5389[16:0], v5390[24:0], v6276[24:0]); // 5.0
    wire [25:0] v6277; shift_adder #(24, 25, 1, 1, 26, 0, 0) op_6277 (v5391[23:0], v4540[24:0], v6277[25:0]); // 5.0
    wire [28:0] v6278; shift_adder #(20, 28, 1, 1, 29, -7, 0) op_6278 (v5392[19:0], v5393[27:0], v6278[28:0]); // 5.0
    wire [28:0] v6279; shift_adder #(26, 24, 1, 1, 29, 4, 0) op_6279 (v5394[25:0], v5395[23:0], v6279[28:0]); // 5.0
    wire [32:0] v6280; shift_adder #(25, 32, 1, 1, 33, -6, 0) op_6280 (v5396[24:0], v5397[31:0], v6280[32:0]); // 5.0
    wire [37:0] v6281; shift_adder #(35, 37, 1, 1, 38, -2, 0) op_6281 (v5398[34:0], v5399[36:0], v6281[37:0]); // 5.0
    wire [19:0] v6282; shift_adder #(18, 14, 1, 1, 20, 5, 0) op_6282 (v5400[17:0], v5401[13:0], v6282[19:0]); // 5.0
    wire [36:0] v6283; shift_adder #(33, 36, 1, 1, 37, -3, 0) op_6283 (v5403[32:0], v5404[35:0], v6283[36:0]); // 5.0
    wire [37:0] v6284; shift_adder #(38, 14, 1, 1, 38, 2, 1) op_6284 (v5405[37:0], v5406[13:0], v6284[37:0]); // 5.0
    wire [21:0] v6285; shift_adder #(21, 19, 1, 1, 22, 2, 0) op_6285 (v5407[20:0], v4484[18:0], v6285[21:0]); // 5.0
    wire [22:0] v6286; shift_adder #(22, 19, 1, 1, 23, 2, 0) op_6286 (v5408[21:0], v5409[18:0], v6286[22:0]); // 5.0
    wire [22:0] v6287; shift_adder #(21, 21, 1, 1, 23, 1, 0) op_6287 (v5410[20:0], v5411[20:0], v6287[22:0]); // 5.0
    wire [18:0] v6288; shift_adder #(18, 17, 1, 1, 19, -1, 0) op_6288 (v5412[17:0], v5413[16:0], v6288[18:0]); // 5.0
    wire [35:0] v6289; shift_adder #(35, 18, 1, 1, 36, 17, 0) op_6289 (v4548[34:0], v5414[17:0], v6289[35:0]); // 5.0
    wire [19:0] v6290; shift_adder #(19, 18, 1, 1, 20, 1, 0) op_6290 (v5415[18:0], v5416[17:0], v6290[19:0]); // 5.0
    wire [34:0] v6291; shift_adder #(34, 22, 1, 1, 35, 11, 0) op_6291 (v5417[33:0], v5418[21:0], v6291[34:0]); // 5.0
    wire [29:0] v6292; shift_adder #(28, 28, 1, 1, 30, -1, 0) op_6292 (v5419[27:0], v5420[27:0], v6292[29:0]); // 5.0
    wire [29:0] v6293; shift_adder #(28, 24, 1, 1, 30, 5, 0) op_6293 (v5421[27:0], v4742[23:0], v6293[29:0]); // 5.0
    wire [21:0] v6294; shift_adder #(19, 19, 1, 1, 22, -3, 0) op_6294 (v5422[18:0], v5423[18:0], v6294[21:0]); // 5.0
    wire [23:0] v6295; shift_adder #(24, 21, 1, 1, 24, 1, 0) op_6295 (v5424[23:0], v5425[20:0], v6295[23:0]); // 5.0
    wire [26:0] v6296; shift_adder #(27, 24, 1, 1, 27, 1, 0) op_6296 (v5426[26:0], v5427[23:0], v6296[26:0]); // 5.0
    wire [24:0] v6297; shift_adder #(23, 15, 1, 1, 25, 9, 0) op_6297 (v5428[22:0], v5429[14:0], v6297[24:0]); // 5.0
    wire [27:0] v6298; shift_adder #(27, 27, 1, 1, 28, 1, 0) op_6298 (v5430[26:0], v5431[26:0], v6298[27:0]); // 5.0
    wire [25:0] v6299; shift_adder #(25, 18, 1, 1, 26, 7, 0) op_6299 (v5432[24:0], v4922[17:0], v6299[25:0]); // 5.0
    wire [22:0] v6300; shift_adder #(18, 23, 1, 1, 23, -3, 0) op_6300 (v5433[17:0], v5434[22:0], v6300[22:0]); // 5.0
    wire [29:0] v6301; shift_adder #(27, 29, 1, 1, 30, -2, 0) op_6301 (v5435[26:0], v5436[28:0], v6301[29:0]); // 5.0
    wire [28:0] v6302; shift_adder #(28, 20, 1, 1, 29, 8, 0) op_6302 (v4989[27:0], v5437[19:0], v6302[28:0]); // 5.0
    wire [33:0] v6303; shift_adder #(33, 32, 1, 1, 34, 2, 0) op_6303 (v4958[32:0], v5438[31:0], v6303[33:0]); // 5.0
    wire [31:0] v6304; shift_adder #(25, 31, 1, 1, 32, -5, 0) op_6304 (v5439[24:0], v5440[30:0], v6304[31:0]); // 5.0
    wire [41:0] v6305; shift_adder #(39, 41, 1, 1, 42, -2, 0) op_6305 (v5441[38:0], v5442[40:0], v6305[41:0]); // 5.0
    wire [18:0] v6306; shift_adder #(17, 16, 1, 1, 19, -2, 0) op_6306 (v5443[16:0], v5444[15:0], v6306[18:0]); // 5.0
    wire [18:0] v6307; shift_adder #(19, 18, 1, 1, 19, 0, 0) op_6307 (v5445[18:0], v5446[17:0], v6307[18:0]); // 5.0
    wire [20:0] v6308; shift_adder #(19, 21, 1, 1, 21, -1, 0) op_6308 (v5447[18:0], v5204[20:0], v6308[20:0]); // 5.0
    wire [19:0] v6309; shift_adder #(17, 18, 1, 1, 20, 2, 0) op_6309 (v5448[16:0], v5449[17:0], v6309[19:0]); // 5.0
    wire [36:0] v6310; shift_adder #(35, 34, 1, 1, 37, 2, 0) op_6310 (v5451[34:0], v5452[33:0], v6310[36:0]); // 5.0
    wire [35:0] v6311; shift_adder #(25, 35, 1, 1, 36, -10, 0) op_6311 (v5453[24:0], v5454[34:0], v6311[35:0]); // 5.0
    wire [32:0] v6312; shift_adder #(33, 20, 1, 1, 33, 12, 0) op_6312 (v5455[32:0], v4724[19:0], v6312[32:0]); // 5.0
    wire [28:0] v6313; shift_adder #(16, 28, 1, 1, 29, -12, 0) op_6313 (v5456[15:0], v5457[27:0], v6313[28:0]); // 5.0
    wire [30:0] v6314; shift_adder #(30, 26, 1, 1, 31, 5, 0) op_6314 (v5458[29:0], v5459[25:0], v6314[30:0]); // 5.0
    wire [31:0] v6315; shift_adder #(31, 28, 1, 1, 32, 2, 0) op_6315 (v5460[30:0], v5461[27:0], v6315[31:0]); // 5.0
    wire [28:0] v6316; shift_adder #(27, 19, 1, 1, 29, 9, 0) op_6316 (v5178[26:0], v5462[18:0], v6316[28:0]); // 5.0
    wire [25:0] v6317; shift_adder #(17, 22, 1, 1, 26, -9, 0) op_6317 (v4794[16:0], v5463[21:0], v6317[25:0]); // 5.0
    wire [22:0] v6318; shift_adder #(16, 21, 1, 1, 23, -6, 0) op_6318 (v5464[15:0], v5465[20:0], v6318[22:0]); // 5.0
    wire [18:0] v6319; shift_adder #(16, 19, 1, 1, 19, -1, 0) op_6319 (v5466[15:0], v5467[18:0], v6319[18:0]); // 5.0
    wire [23:0] v6320; shift_adder #(21, 17, 1, 1, 24, 7, 0) op_6320 (v5468[20:0], v5469[16:0], v6320[23:0]); // 5.0
    wire [24:0] v6321; shift_adder #(21, 25, 1, 1, 25, -1, 0) op_6321 (v5470[20:0], v5471[24:0], v6321[24:0]); // 5.0
    wire [33:0] v6322; shift_adder #(21, 33, 1, 1, 34, -11, 0) op_6322 (v5472[20:0], v5473[32:0], v6322[33:0]); // 5.0
    wire [27:0] v6323; shift_adder #(26, 16, 1, 1, 28, 11, 0) op_6323 (v5474[25:0], v5475[15:0], v6323[27:0]); // 5.0
    wire [31:0] v6324; shift_adder #(26, 30, 1, 1, 32, -5, 0) op_6324 (v5476[25:0], v5477[29:0], v6324[31:0]); // 5.0
    wire [34:0] v6325; shift_adder #(24, 34, 1, 1, 35, -9, 0) op_6325 (v5478[23:0], v5479[33:0], v6325[34:0]); // 5.0
    wire [28:0] v6326; shift_adder #(28, 19, 1, 1, 29, 8, 0) op_6326 (v5480[27:0], v5229[18:0], v6326[28:0]); // 5.0
    wire [38:0] v6327; shift_adder #(37, 38, 1, 1, 39, -2, 0) op_6327 (v5481[36:0], v5482[37:0], v6327[38:0]); // 5.0
    wire [36:0] v6328; shift_adder #(37, 18, 1, 1, 37, 0, 1) op_6328 (v5483[36:0], v5484[17:0], v6328[36:0]); // 5.0
    wire [36:0] v6329; shift_adder #(17, 37, 1, 1, 37, -18, 0) op_6329 (v5485[16:0], v5486[36:0], v6329[36:0]); // 5.0
    wire [21:0] v6330; shift_adder #(19, 20, 1, 1, 22, -2, 0) op_6330 (v5487[18:0], v5488[19:0], v6330[21:0]); // 5.0
    wire [18:0] v6331; shift_adder #(18, 17, 1, 1, 19, -1, 0) op_6331 (v5489[17:0], v5490[16:0], v6331[18:0]); // 5.0
    wire [31:0] v6332; shift_adder #(17, 31, 1, 1, 32, -14, 0) op_6332 (v5491[16:0], v5492[30:0], v6332[31:0]); // 5.0
    wire [27:0] v6333; shift_adder #(27, 27, 1, 1, 28, 0, 0) op_6333 (v5493[26:0], v5494[26:0], v6333[27:0]); // 5.0
    wire [28:0] v6334; shift_adder #(19, 27, 1, 1, 29, -9, 0) op_6334 (v5495[18:0], v4749[26:0], v6334[28:0]); // 5.0
    wire [28:0] v6335; shift_adder #(28, 27, 1, 1, 29, 1, 0) op_6335 (v4455[27:0], v5496[26:0], v6335[28:0]); // 5.0
    wire [27:0] v6336; shift_adder #(27, 16, 1, 1, 28, 11, 0) op_6336 (v5497[26:0], v5498[15:0], v6336[27:0]); // 5.0
    wire [24:0] v6337; shift_adder #(24, 22, 1, 1, 25, 2, 0) op_6337 (v5499[23:0], v5500[21:0], v6337[24:0]); // 5.0
    wire [21:0] v6338; shift_adder #(21, 21, 1, 1, 22, 0, 0) op_6338 (v5501[20:0], v5502[20:0], v6338[21:0]); // 5.0
    wire [23:0] v6339; shift_adder #(19, 18, 1, 1, 24, 6, 0) op_6339 (v5503[18:0], v5504[17:0], v6339[23:0]); // 5.0
    wire [22:0] v6340; shift_adder #(17, 22, 1, 1, 23, -4, 0) op_6340 (v5505[16:0], v5506[21:0], v6340[22:0]); // 5.0
    wire [20:0] v6341; shift_adder #(19, 18, 1, 1, 21, 2, 0) op_6341 (v5507[18:0], v5508[17:0], v6341[20:0]); // 5.0
    wire [24:0] v6342; shift_adder #(22, 24, 1, 1, 25, -2, 0) op_6342 (v5509[21:0], v5510[23:0], v6342[24:0]); // 5.0
    wire [26:0] v6343; shift_adder #(24, 26, 1, 1, 27, -2, 0) op_6343 (v5511[23:0], v5276[25:0], v6343[26:0]); // 5.0
    wire [32:0] v6344; shift_adder #(25, 32, 1, 1, 33, -7, 0) op_6344 (v5512[24:0], v5513[31:0], v6344[32:0]); // 5.0
    wire [34:0] v6345; shift_adder #(21, 34, 1, 1, 35, -12, 0) op_6345 (v5514[20:0], v5515[33:0], v6345[34:0]); // 5.0
    wire [38:0] v6346; shift_adder #(39, 17, 1, 1, 39, 3, 1) op_6346 (v5516[38:0], v5517[16:0], v6346[38:0]); // 5.0
    wire [25:0] v6347; shift_adder #(21, 23, 1, 1, 26, -4, 0) op_6347 (v5518[20:0], v5519[22:0], v6347[25:0]); // 5.0
    wire [22:0] v6348; shift_adder #(20, 19, 1, 1, 23, -3, 0) op_6348 (v5520[19:0], v5521[18:0], v6348[22:0]); // 5.0
    wire [33:0] v6349; shift_adder #(32, 16, 1, 1, 34, 18, 0) op_6349 (v5522[31:0], v5523[15:0], v6349[33:0]); // 5.0
    wire [37:0] v6350; shift_adder #(16, 14, 1, 1, 38, 24, 1) op_6350 (v5524[15:0], v4152[13:0], v6350[37:0]); // 5.0
    wire [32:0] v6351; shift_adder #(21, 32, 1, 1, 33, -11, 0) op_6351 (v5525[20:0], v5088[31:0], v6351[32:0]); // 5.0
    wire [40:0] v6352; shift_adder #(40, 36, 1, 1, 41, 4, 0) op_6352 (v5526[39:0], v5527[35:0], v6352[40:0]); // 5.0
    wire [32:0] v6353; shift_adder #(24, 32, 1, 1, 33, -7, 0) op_6353 (v5528[23:0], v5529[31:0], v6353[32:0]); // 5.0
    wire [28:0] v6354; shift_adder #(28, 27, 1, 1, 29, -1, 0) op_6354 (v5530[27:0], v5531[26:0], v6354[28:0]); // 5.0
    wire [33:0] v6355; shift_adder #(33, 33, 1, 1, 34, 0, 0) op_6355 (v5532[32:0], v4596[32:0], v6355[33:0]); // 5.0
    wire [30:0] v6356; shift_adder #(31, 16, 1, 1, 31, 12, 0) op_6356 (v5533[30:0], v5534[15:0], v6356[30:0]); // 5.0
    wire [32:0] v6357; shift_adder #(32, 25, 1, 1, 33, 7, 0) op_6357 (v5034[31:0], v5535[24:0], v6357[32:0]); // 5.0
    wire [29:0] v6358; shift_adder #(29, 19, 1, 1, 30, 10, 0) op_6358 (v5536[28:0], v5537[18:0], v6358[29:0]); // 5.0
    wire [28:0] v6359; shift_adder #(24, 26, 1, 1, 29, -5, 0) op_6359 (v5538[23:0], v5539[25:0], v6359[28:0]); // 5.0
    wire [23:0] v6360; shift_adder #(24, 18, 1, 1, 24, 4, 0) op_6360 (v5011[23:0], v5540[17:0], v6360[23:0]); // 5.0
    wire [24:0] v6361; shift_adder #(23, 23, 1, 1, 25, 1, 0) op_6361 (v5541[22:0], v4545[22:0], v6361[24:0]); // 5.0
    wire [25:0] v6362; shift_adder #(24, 23, 1, 1, 26, 2, 0) op_6362 (v5542[23:0], v5543[22:0], v6362[25:0]); // 5.0
    wire [30:0] v6363; shift_adder #(29, 29, 1, 1, 31, 2, 0) op_6363 (v5544[28:0], v5545[28:0], v6363[30:0]); // 5.0
    wire [19:0] v6364; shift_adder #(19, 18, 1, 1, 20, 1, 0) op_6364 (v4861[18:0], v5546[17:0], v6364[19:0]); // 5.0
    wire [28:0] v6365; shift_adder #(19, 27, 1, 1, 29, -10, 0) op_6365 (v5547[18:0], v5548[26:0], v6365[28:0]); // 5.0
    wire [27:0] v6366; shift_adder #(27, 25, 1, 1, 28, 1, 0) op_6366 (v5549[26:0], v5550[24:0], v6366[27:0]); // 5.0
    wire [25:0] v6367; shift_adder #(20, 25, 1, 1, 26, -5, 0) op_6367 (v4494[19:0], v5551[24:0], v6367[25:0]); // 5.0
    wire [28:0] v6368; shift_adder #(29, 27, 1, 1, 29, 0, 0) op_6368 (v5552[28:0], v5553[26:0], v6368[28:0]); // 5.0
    wire [31:0] v6369; shift_adder #(30, 23, 1, 1, 32, 8, 0) op_6369 (v5554[29:0], v5555[22:0], v6369[31:0]); // 5.0
    wire [29:0] v6370; shift_adder #(27, 20, 1, 1, 30, 9, 0) op_6370 (v5556[26:0], v5557[19:0], v6370[29:0]); // 5.0
    wire [33:0] v6371; shift_adder #(29, 33, 1, 1, 34, -3, 0) op_6371 (v4800[28:0], v5558[32:0], v6371[33:0]); // 5.0
    wire [35:0] v6372; shift_adder #(28, 36, 1, 1, 36, -6, 0) op_6372 (v5207[27:0], v5559[35:0], v6372[35:0]); // 5.0
    wire [23:0] v6373; shift_adder #(20, 21, 1, 1, 24, 3, 0) op_6373 (v5560[19:0], v5561[20:0], v6373[23:0]); // 5.0
    wire [32:0] v6374; shift_adder #(29, 32, 1, 1, 33, -3, 0) op_6374 (v5563[28:0], v5513[31:0], v6374[32:0]); // 5.0
    wire [40:0] v6375; shift_adder #(40, 18, 1, 1, 41, 22, 0) op_6375 (v5564[39:0], v5565[17:0], v6375[40:0]); // 5.0
    wire [39:0] v6376; shift_adder #(39, 15, 1, 1, 40, 24, 0) op_6376 (v5566[38:0], v5567[14:0], v6376[39:0]); // 5.0
    wire [17:0] v6377; shift_adder #(17, 15, 1, 1, 18, 1, 0) op_6377 (v4547[16:0], v5568[14:0], v6377[17:0]); // 5.0
    wire [22:0] v6378; shift_adder #(22, 22, 1, 1, 23, 1, 0) op_6378 (v5569[21:0], v4865[21:0], v6378[22:0]); // 5.0
    wire [25:0] v6379; shift_adder #(26, 23, 1, 1, 26, 1, 0) op_6379 (v5570[25:0], v5571[22:0], v6379[25:0]); // 5.0
    wire [22:0] v6380; shift_adder #(20, 20, 1, 1, 23, -2, 0) op_6380 (v5572[19:0], v5573[19:0], v6380[22:0]); // 5.0
    wire [17:0] v6381; shift_adder #(16, 16, 1, 1, 18, -2, 0) op_6381 (v5574[15:0], v5575[15:0], v6381[17:0]); // 5.0
    wire [20:0] v6382; shift_adder #(17, 20, 1, 1, 21, -1, 0) op_6382 (v5576[16:0], v5577[19:0], v6382[20:0]); // 5.0
    wire [22:0] v6383; shift_adder #(22, 21, 1, 1, 23, 1, 0) op_6383 (v5578[21:0], v5579[20:0], v6383[22:0]); // 5.0
    wire [23:0] v6384; shift_adder #(22, 23, 1, 1, 24, -1, 0) op_6384 (v5580[21:0], v5581[22:0], v6384[23:0]); // 5.0
    wire [25:0] v6385; shift_adder #(24, 21, 1, 1, 26, 4, 0) op_6385 (v5582[23:0], v5583[20:0], v6385[25:0]); // 5.0
    wire [29:0] v6386; shift_adder #(28, 29, 1, 1, 30, 0, 0) op_6386 (v5584[27:0], v5585[28:0], v6386[29:0]); // 5.0
    wire [30:0] v6387; shift_adder #(28, 19, 1, 1, 31, 12, 0) op_6387 (v4815[27:0], v5586[18:0], v6387[30:0]); // 5.0
    wire [28:0] v6388; shift_adder #(27, 27, 1, 1, 29, 1, 0) op_6388 (v5587[26:0], v4842[26:0], v6388[28:0]); // 5.0
    wire [31:0] v6389; shift_adder #(28, 31, 1, 1, 32, -3, 0) op_6389 (v5588[27:0], v5589[30:0], v6389[31:0]); // 5.0
    wire [36:0] v6390; shift_adder #(16, 17, 1, 1, 37, 20, 1) op_6390 (v5590[15:0], v4239[16:0], v6390[36:0]); // 5.0
    wire [22:0] v6391; shift_adder #(21, 19, 1, 1, 23, 4, 0) op_6391 (v5591[20:0], v5592[18:0], v6391[22:0]); // 5.0
    wire [36:0] v6392; shift_adder #(25, 36, 1, 1, 37, -11, 0) op_6392 (v5593[24:0], v5594[35:0], v6392[36:0]); // 5.0
    wire [38:0] v6393; shift_adder #(38, 29, 1, 1, 39, 9, 0) op_6393 (v5595[37:0], v5596[28:0], v6393[38:0]); // 5.0
    wire [38:0] v6394; shift_adder #(16, 15, 1, 1, 39, -23, 1) op_6394 (v5597[15:0], v5598[14:0], v6394[38:0]); // 5.0
    wire [20:0] v6395; shift_adder #(16, 16, 1, 1, 21, -4, 0) op_6395 (v5599[15:0], v5600[15:0], v6395[20:0]); // 5.0
    wire [34:0] v6396; shift_adder #(34, 32, 1, 1, 35, 2, 0) op_6396 (v5601[33:0], v5602[31:0], v6396[34:0]); // 5.0
    wire [28:0] v6397; shift_adder #(22, 28, 1, 1, 29, -5, 0) op_6397 (v5603[21:0], v5604[27:0], v6397[28:0]); // 5.0
    wire [27:0] v6398; shift_adder #(27, 26, 1, 1, 28, -1, 0) op_6398 (v5112[26:0], v5605[25:0], v6398[27:0]); // 5.0
    wire [27:0] v6399; shift_adder #(27, 26, 1, 1, 28, 0, 0) op_6399 (v5606[26:0], v5607[25:0], v6399[27:0]); // 5.0
    wire [22:0] v6400; shift_adder #(23, 17, 1, 1, 23, 5, 0) op_6400 (v5608[22:0], v5609[16:0], v6400[22:0]); // 5.0
    wire [26:0] v6401; shift_adder #(26, 21, 1, 1, 27, 5, 0) op_6401 (v5610[25:0], v5611[20:0], v6401[26:0]); // 5.0
    wire [24:0] v6402; shift_adder #(23, 24, 1, 1, 25, -2, 0) op_6402 (v5612[22:0], v5613[23:0], v6402[24:0]); // 5.0
    wire [20:0] v6403; shift_adder #(20, 18, 1, 1, 21, 1, 0) op_6403 (v5614[19:0], v4901[17:0], v6403[20:0]); // 5.0
    wire [22:0] v6404; shift_adder #(20, 22, 1, 1, 23, 0, 0) op_6404 (v5615[19:0], v5616[21:0], v6404[22:0]); // 5.0
    wire [29:0] v6405; shift_adder #(26, 30, 1, 1, 30, -2, 0) op_6405 (v5617[25:0], v5618[29:0], v6405[29:0]); // 5.0
    wire [32:0] v6406; shift_adder #(30, 29, 1, 1, 33, 3, 0) op_6406 (v5619[29:0], v5620[28:0], v6406[32:0]); // 5.0
    wire [24:0] v6407; shift_adder #(23, 23, 1, 1, 25, 2, 0) op_6407 (v5621[22:0], v5622[22:0], v6407[24:0]); // 5.0
    wire [25:0] v6408; shift_adder #(20, 26, 1, 1, 26, -3, 0) op_6408 (v5623[19:0], v5624[25:0], v6408[25:0]); // 5.0
    wire [24:0] v6409; shift_adder #(24, 19, 1, 1, 25, 5, 0) op_6409 (v5625[23:0], v5626[18:0], v6409[24:0]); // 5.0
    wire [23:0] v6410; shift_adder #(23, 18, 1, 1, 24, 4, 0) op_6410 (v5627[22:0], v5628[17:0], v6410[23:0]); // 5.0
    wire [37:0] v6411; shift_adder #(15, 19, 1, 1, 38, 19, 1) op_6411 (v5629[14:0], v4286[18:0], v6411[37:0]); // 5.0
    wire [39:0] v6412; shift_adder #(39, 21, 1, 1, 40, 19, 0) op_6412 (v5630[38:0], v5631[20:0], v6412[39:0]); // 5.0
    wire [19:0] v6413; shift_adder #(19, 17, 1, 1, 20, 0, 0) op_6413 (v5632[18:0], v4458[16:0], v6413[19:0]); // 5.0
    wire [21:0] v6414; shift_adder #(21, 18, 1, 1, 22, 2, 0) op_6414 (v5633[20:0], v5634[17:0], v6414[21:0]); // 5.0
    wire [29:0] v6415; shift_adder #(28, 29, 1, 1, 30, -1, 0) op_6415 (v5457[27:0], v4613[28:0], v6415[29:0]); // 5.0
    wire [41:0] v6416; shift_adder #(42, 19, 1, 1, 42, 3, 1) op_6416 (v5635[41:0], v5636[18:0], v6416[41:0]); // 5.0
    wire [18:0] v6417; shift_adder #(16, 17, 1, 1, 19, 2, 0) op_6417 (v5637[15:0], v5638[16:0], v6417[18:0]); // 5.0
    wire [32:0] v6418; shift_adder #(27, 33, 1, 1, 33, -5, 0) op_6418 (v4457[26:0], v5640[32:0], v6418[32:0]); // 5.0
    wire [32:0] v6419; shift_adder #(31, 19, 1, 1, 33, 14, 0) op_6419 (v5589[30:0], v5641[18:0], v6419[32:0]); // 5.0
    wire [25:0] v6420; shift_adder #(23, 24, 1, 1, 26, -2, 0) op_6420 (v4482[22:0], v5642[23:0], v6420[25:0]); // 5.0
    wire [30:0] v6421; shift_adder #(30, 29, 1, 1, 31, 2, 0) op_6421 (v5643[29:0], v5644[28:0], v6421[30:0]); // 5.0
    wire [29:0] v6422; shift_adder #(23, 29, 1, 1, 30, -6, 0) op_6422 (v5645[22:0], v5100[28:0], v6422[29:0]); // 5.0
    wire [30:0] v6423; shift_adder #(30, 28, 1, 1, 31, 1, 0) op_6423 (v5646[29:0], v5647[27:0], v6423[30:0]); // 5.0
    wire [27:0] v6424; shift_adder #(25, 27, 1, 1, 28, -2, 0) op_6424 (v5648[24:0], v5649[26:0], v6424[27:0]); // 5.0
    wire [21:0] v6425; shift_adder #(18, 19, 1, 1, 22, -3, 0) op_6425 (v5650[17:0], v5651[18:0], v6425[21:0]); // 5.0
    wire [19:0] v6426; shift_adder #(17, 18, 1, 1, 20, 2, 0) op_6426 (v5652[16:0], v5653[17:0], v6426[19:0]); // 5.0
    wire [19:0] v6427; shift_adder #(18, 16, 1, 1, 20, 3, 0) op_6427 (v5654[17:0], v5655[15:0], v6427[19:0]); // 5.0
    wire [24:0] v6428; shift_adder #(20, 16, 1, 1, 25, 9, 0) op_6428 (v5656[19:0], v5657[15:0], v6428[24:0]); // 5.0
    wire [24:0] v6429; shift_adder #(22, 25, 1, 1, 25, -1, 0) op_6429 (v5658[21:0], v5659[24:0], v6429[24:0]); // 5.0
    wire [31:0] v6430; shift_adder #(31, 23, 1, 1, 32, 8, 0) op_6430 (v5660[30:0], v5661[22:0], v6430[31:0]); // 5.0
    wire [32:0] v6431; shift_adder #(31, 30, 1, 1, 33, 2, 0) op_6431 (v5662[30:0], v5663[29:0], v6431[32:0]); // 5.0
    wire [29:0] v6432; shift_adder #(28, 16, 1, 1, 30, 13, 0) op_6432 (v4662[27:0], v5664[15:0], v6432[29:0]); // 5.0
    wire [31:0] v6433; shift_adder #(28, 31, 1, 1, 32, -2, 0) op_6433 (v5665[27:0], v5666[30:0], v6433[31:0]); // 5.0
    wire [32:0] v6434; shift_adder #(32, 26, 1, 1, 33, 7, 0) op_6434 (v5667[31:0], v4947[25:0], v6434[32:0]); // 5.0
    wire [25:0] v6435; shift_adder #(24, 20, 1, 1, 26, 5, 0) op_6435 (v5668[23:0], v5669[19:0], v6435[25:0]); // 5.0
    wire [32:0] v6436; shift_adder #(32, 27, 1, 1, 33, 5, 0) op_6436 (v5670[31:0], v5167[26:0], v6436[32:0]); // 5.0
    wire [30:0] v6437; shift_adder #(26, 30, 1, 1, 31, -4, 0) op_6437 (v5671[25:0], v5672[29:0], v6437[30:0]); // 5.0
    wire [30:0] v6438; shift_adder #(29, 30, 1, 1, 31, -1, 0) op_6438 (v5673[28:0], v5674[29:0], v6438[30:0]); // 5.0
    wire [38:0] v6439; shift_adder #(21, 39, 1, 1, 39, -17, 0) op_6439 (v5675[20:0], v5676[38:0], v6439[38:0]); // 5.0
    wire [31:0] v6440; shift_adder #(31, 24, 1, 1, 32, 6, 0) op_6440 (v5677[30:0], v5678[23:0], v6440[31:0]); // 5.0
    wire [30:0] v6441; shift_adder #(18, 29, 1, 1, 31, -13, 0) op_6441 (v5679[17:0], v5680[28:0], v6441[30:0]); // 5.0
    wire [25:0] v6442; shift_adder #(23, 25, 1, 1, 26, -2, 0) op_6442 (v5681[22:0], v5132[24:0], v6442[25:0]); // 5.0
    wire [29:0] v6443; shift_adder #(29, 28, 1, 1, 30, 0, 0) op_6443 (v5682[28:0], v5683[27:0], v6443[29:0]); // 5.0
    wire [22:0] v6444; shift_adder #(23, 21, 1, 1, 23, 0, 0) op_6444 (v5684[22:0], v5685[20:0], v6444[22:0]); // 5.0
    wire [23:0] v6445; shift_adder #(23, 18, 1, 1, 24, 3, 0) op_6445 (v5686[22:0], v5687[17:0], v6445[23:0]); // 5.0
    wire [19:0] v6446; shift_adder #(19, 18, 1, 1, 20, -1, 0) op_6446 (v5688[18:0], v5689[17:0], v6446[19:0]); // 5.0
    wire [16:0] v6447; shift_adder #(17, 16, 1, 1, 17, 0, 0) op_6447 (v5690[16:0], v5691[15:0], v6447[16:0]); // 5.0
    wire [20:0] v6448; shift_adder #(18, 19, 1, 1, 21, 1, 0) op_6448 (v5692[17:0], v5693[18:0], v6448[20:0]); // 5.0
    wire [22:0] v6449; shift_adder #(22, 20, 1, 1, 23, 3, 0) op_6449 (v5694[21:0], v5695[19:0], v6449[22:0]); // 5.0
    wire [24:0] v6450; shift_adder #(23, 25, 1, 1, 25, 0, 0) op_6450 (v5696[22:0], v5697[24:0], v6450[24:0]); // 5.0
    wire [23:0] v6451; shift_adder #(22, 23, 1, 1, 24, 0, 0) op_6451 (v5698[21:0], v5699[22:0], v6451[23:0]); // 5.0
    wire [26:0] v6452; shift_adder #(25, 24, 1, 1, 27, 2, 0) op_6452 (v5700[24:0], v5701[23:0], v6452[26:0]); // 5.0
    wire [31:0] v6453; shift_adder #(26, 32, 1, 1, 32, -5, 0) op_6453 (v5702[25:0], v5703[31:0], v6453[31:0]); // 5.0
    wire [26:0] v6454; shift_adder #(26, 17, 1, 1, 27, 9, 0) op_6454 (v5215[25:0], v5704[16:0], v6454[26:0]); // 5.0
    wire [30:0] v6455; shift_adder #(29, 25, 1, 1, 31, 6, 0) op_6455 (v5705[28:0], v5706[24:0], v6455[30:0]); // 5.0
    wire [24:0] v6456; shift_adder #(23, 21, 1, 1, 25, 3, 0) op_6456 (v5707[22:0], v5708[20:0], v6456[24:0]); // 5.0
    wire [32:0] v6457; shift_adder #(28, 32, 1, 1, 33, -3, 0) op_6457 (v5709[27:0], v5710[31:0], v6457[32:0]); // 5.0
    wire [33:0] v6458; shift_adder #(27, 34, 1, 1, 34, -5, 0) op_6458 (v5711[26:0], v5712[33:0], v6458[33:0]); // 5.0
    wire [34:0] v6459; shift_adder #(33, 28, 1, 1, 35, 6, 0) op_6459 (v5713[32:0], v5714[27:0], v6459[34:0]); // 5.0
    wire [40:0] v6460; shift_adder #(40, 25, 1, 1, 41, 16, 0) op_6460 (v5715[39:0], v5716[24:0], v6460[40:0]); // 5.0
    wire [38:0] v6461; shift_adder #(37, 38, 1, 1, 39, 0, 0) op_6461 (v5717[36:0], v5718[37:0], v6461[38:0]); // 5.0
    wire [27:0] v6462; shift_adder #(15, 28, 1, 1, 28, -11, 0) op_6462 (v5719[14:0], v5720[27:0], v6462[27:0]); // 5.0
    wire [33:0] v6463; shift_adder #(27, 31, 1, 1, 34, -7, 0) op_6463 (v5426[26:0], v5721[30:0], v6463[33:0]); // 5.0
    wire [26:0] v6464; shift_adder #(21, 26, 1, 1, 27, -6, 0) op_6464 (v5722[20:0], v5723[25:0], v6464[26:0]); // 5.0
    wire [28:0] v6465; shift_adder #(28, 17, 1, 1, 29, 10, 0) op_6465 (v5724[27:0], v4721[16:0], v6465[28:0]); // 5.0
    wire [28:0] v6466; shift_adder #(21, 27, 1, 1, 29, -7, 0) op_6466 (v5725[20:0], v4986[26:0], v6466[28:0]); // 5.0
    wire [25:0] v6467; shift_adder #(22, 25, 1, 1, 26, -4, 0) op_6467 (v5726[21:0], v5727[24:0], v6467[25:0]); // 5.0
    wire [19:0] v6468; shift_adder #(18, 19, 1, 1, 20, -1, 0) op_6468 (v5728[17:0], v5729[18:0], v6468[19:0]); // 5.0
    wire [21:0] v6469; shift_adder #(22, 17, 1, 1, 22, 2, 0) op_6469 (v5730[21:0], v5731[16:0], v6469[21:0]); // 5.0
    wire [29:0] v6470; shift_adder #(24, 30, 1, 1, 30, -2, 0) op_6470 (v5732[23:0], v5733[29:0], v6470[29:0]); // 5.0
    wire [29:0] v6471; shift_adder #(18, 29, 1, 1, 30, -10, 0) op_6471 (v5650[17:0], v5734[28:0], v6471[29:0]); // 5.0
    wire [26:0] v6472; shift_adder #(25, 26, 1, 1, 27, 1, 0) op_6472 (v5735[24:0], v5736[25:0], v6472[26:0]); // 5.0
    wire [23:0] v6473; shift_adder #(22, 18, 1, 1, 24, 6, 0) op_6473 (v5737[21:0], v5738[17:0], v6473[23:0]); // 5.0
    wire [22:0] v6474; shift_adder #(15, 23, 1, 1, 23, -6, 0) op_6474 (v5739[14:0], v5740[22:0], v6474[22:0]); // 5.0
    wire [30:0] v6475; shift_adder #(30, 23, 1, 1, 31, 7, 0) op_6475 (v5741[29:0], v5742[22:0], v6475[30:0]); // 5.0
    wire [33:0] v6476; shift_adder #(30, 33, 1, 1, 34, -1, 0) op_6476 (v5743[29:0], v5744[32:0], v6476[33:0]); // 5.0
    wire [38:0] v6477; shift_adder #(37, 17, 1, 1, 39, -2, 1) op_6477 (v5745[36:0], v5746[16:0], v6477[38:0]); // 5.0
    wire [20:0] v6478; shift_adder #(18, 20, 1, 1, 21, -3, 0) op_6478 (v5747[17:0], v5748[19:0], v6478[20:0]); // 5.0
    wire [23:0] v6479; shift_adder #(22, 17, 1, 1, 24, 6, 0) op_6479 (v5749[21:0], v5750[16:0], v6479[23:0]); // 5.0
    wire [36:0] v6480; shift_adder #(18, 18, 1, 1, 37, 19, 1) op_6480 (v5751[17:0], v4427[17:0], v6480[36:0]); // 5.0
    wire [27:0] v6481; shift_adder #(20, 28, 1, 1, 28, -7, 0) op_6481 (v5752[19:0], v5753[27:0], v6481[27:0]); // 5.0
    wire [37:0] v6482; shift_adder #(37, 36, 1, 1, 38, 0, 0) op_6482 (v5754[36:0], v5755[35:0], v6482[37:0]); // 5.0
    wire [33:0] v6483; shift_adder #(34, 25, 1, 1, 34, 8, 0) op_6483 (v5756[33:0], v5128[24:0], v6483[33:0]); // 5.0
    wire [38:0] v6484; shift_adder #(38, 32, 1, 1, 39, 5, 0) op_6484 (v5757[37:0], v5758[31:0], v6484[38:0]); // 5.0
    wire [26:0] v6485; shift_adder #(26, 25, 1, 1, 27, 0, 0) op_6485 (v5759[25:0], v5760[24:0], v6485[26:0]); // 5.0
    wire [28:0] v6486; shift_adder #(19, 28, 1, 1, 29, -10, 0) op_6486 (v5761[18:0], v5762[27:0], v6486[28:0]); // 5.0
    wire [34:0] v6487; shift_adder #(26, 32, 1, 1, 35, -8, 0) op_6487 (v5763[25:0], v5764[31:0], v6487[34:0]); // 5.0
    wire [29:0] v6488; shift_adder #(15, 30, 1, 1, 30, -14, 0) op_6488 (v5765[14:0], v5766[29:0], v6488[29:0]); // 5.0
    wire [24:0] v6489; shift_adder #(25, 17, 1, 1, 25, 6, 0) op_6489 (v5767[24:0], v5768[16:0], v6489[24:0]); // 5.0
    wire [23:0] v6490; shift_adder #(20, 20, 1, 1, 24, -4, 0) op_6490 (v5769[19:0], v5770[19:0], v6490[23:0]); // 5.0
    wire [25:0] v6491; shift_adder #(25, 25, 1, 1, 26, 0, 0) op_6491 (v5771[24:0], v5772[24:0], v6491[25:0]); // 6.0
    wire [29:0] v6492; shift_adder #(26, 30, 1, 1, 30, -2, 0) op_6492 (v5773[25:0], v5774[29:0], v6492[29:0]); // 6.0
    wire [32:0] v6493; shift_adder #(10, 33, 1, 1, 33, -8, 1) op_6493 (v170[9:0], v5775[32:0], v6493[32:0]); // 6.0
    wire [31:0] v6494; shift_adder #(26, 32, 1, 1, 32, -3, 0) op_6494 (v5776[25:0], v5777[31:0], v6494[31:0]); // 6.0
    wire [29:0] v6495; shift_adder #(27, 29, 1, 1, 30, -1, 0) op_6495 (v5778[26:0], v5779[28:0], v6495[29:0]); // 6.0
    wire [32:0] v6496; shift_adder #(33, 26, 1, 1, 33, 3, 0) op_6496 (v5780[32:0], v5781[25:0], v6496[32:0]); // 6.0
    wire [37:0] v6497; shift_adder #(19, 28, 1, 1, 38, 10, 1) op_6497 (v5782[18:0], v4467[27:0], v6497[37:0]); // 6.0
    wire [29:0] v6498; shift_adder #(25, 30, 1, 1, 30, -4, 0) op_6498 (v5783[24:0], v5784[29:0], v6498[29:0]); // 6.0
    wire [25:0] v6499; shift_adder #(24, 23, 1, 1, 26, 3, 0) op_6499 (v5785[23:0], v5786[22:0], v6499[25:0]); // 6.0
    wire [37:0] v6500; shift_adder #(37, 33, 1, 1, 38, 4, 0) op_6500 (v5788[36:0], v5789[32:0], v6500[37:0]); // 6.0
    wire [22:0] v6501; shift_adder #(23, 20, 1, 1, 23, 0, 0) op_6501 (v5790[22:0], v5791[19:0], v6501[22:0]); // 6.0
    wire [32:0] v6502; shift_adder #(32, 27, 1, 1, 33, 4, 0) op_6502 (v5792[31:0], v5793[26:0], v6502[32:0]); // 6.0
    wire [24:0] v6503; shift_adder #(23, 23, 1, 1, 25, -1, 0) op_6503 (v5794[22:0], v5795[22:0], v6503[24:0]); // 6.0
    wire [25:0] v6504; shift_adder #(21, 26, 1, 1, 26, 0, 0) op_6504 (v5796[20:0], v5797[25:0], v6504[25:0]); // 6.0
    wire [29:0] v6505; shift_adder #(27, 30, 1, 1, 30, -1, 0) op_6505 (v5798[26:0], v5799[29:0], v6505[29:0]); // 6.0
    wire [35:0] v6506; shift_adder #(11, 35, 1, 1, 36, -24, 1) op_6506 (v312[10:0], v5800[34:0], v6506[35:0]); // 6.0
    wire [23:0] v6507; shift_adder #(24, 18, 1, 1, 24, 5, 0) op_6507 (v5801[23:0], v5802[17:0], v6507[23:0]); // 6.0
    wire [29:0] v6508; shift_adder #(28, 28, 1, 1, 30, -2, 0) op_6508 (v5803[27:0], v5804[27:0], v6508[29:0]); // 6.0
    wire [33:0] v6509; shift_adder #(30, 33, 1, 1, 34, -2, 0) op_6509 (v5805[29:0], v5806[32:0], v6509[33:0]); // 6.0
    wire [34:0] v6510; shift_adder #(35, 29, 1, 1, 35, 5, 0) op_6510 (v5807[34:0], v5808[28:0], v6510[34:0]); // 6.0
    wire [36:0] v6511; shift_adder #(37, 20, 1, 1, 37, 0, 1) op_6511 (v5809[36:0], v5810[19:0], v6511[36:0]); // 6.0
    wire [24:0] v6512; shift_adder #(24, 22, 1, 1, 25, 2, 0) op_6512 (v5811[23:0], v5812[21:0], v6512[24:0]); // 6.0
    wire [37:0] v6513; shift_adder #(20, 29, 1, 1, 38, 9, 1) op_6513 (v5813[19:0], v4527[28:0], v6513[37:0]); // 6.0
    wire [40:0] v6514; shift_adder #(28, 40, 1, 1, 41, -11, 0) op_6514 (v5814[27:0], v5815[39:0], v6514[40:0]); // 6.0
    wire [29:0] v6515; shift_adder #(29, 25, 1, 1, 30, 3, 0) op_6515 (v5816[28:0], v5817[24:0], v6515[29:0]); // 6.0
    wire [26:0] v6516; shift_adder #(25, 25, 1, 1, 27, -2, 0) op_6516 (v5818[24:0], v5819[24:0], v6516[26:0]); // 6.0
    wire [30:0] v6517; shift_adder #(27, 31, 1, 1, 31, -1, 0) op_6517 (v5820[26:0], v5821[30:0], v6517[30:0]); // 6.0
    wire [30:0] v6518; shift_adder #(29, 26, 1, 1, 31, 4, 0) op_6518 (v5822[28:0], v5823[25:0], v6518[30:0]); // 6.0
    wire [36:0] v6519; shift_adder #(37, 28, 1, 1, 37, 7, 0) op_6519 (v5824[36:0], v5825[27:0], v6519[36:0]); // 6.0
    wire [24:0] v6520; shift_adder #(24, 24, 1, 1, 25, -1, 0) op_6520 (v5826[23:0], v5827[23:0], v6520[24:0]); // 6.0
    wire [32:0] v6521; shift_adder #(32, 28, 1, 1, 33, 3, 0) op_6521 (v5828[31:0], v5829[27:0], v6521[32:0]); // 6.0
    wire [40:0] v6522; shift_adder #(41, 19, 1, 1, 41, 0, 1) op_6522 (v5830[40:0], v5831[18:0], v6522[40:0]); // 6.0
    wire [37:0] v6523; shift_adder #(35, 37, 1, 1, 38, -1, 0) op_6523 (v5832[34:0], v5833[36:0], v6523[37:0]); // 6.0
    wire [31:0] v6524; shift_adder #(24, 30, 1, 1, 32, -8, 0) op_6524 (v5834[23:0], v5835[29:0], v6524[31:0]); // 6.0
    wire [21:0] v6525; shift_adder #(21, 19, 1, 1, 22, -1, 0) op_6525 (v5836[20:0], v5837[18:0], v6525[21:0]); // 6.0
    wire [32:0] v6526; shift_adder #(29, 33, 1, 1, 33, -3, 0) op_6526 (v5838[28:0], v5839[32:0], v6526[32:0]); // 6.0
    wire [34:0] v6527; shift_adder #(34, 29, 1, 1, 35, 5, 0) op_6527 (v5840[33:0], v5841[28:0], v6527[34:0]); // 6.0
    wire [27:0] v6528; shift_adder #(24, 23, 1, 1, 28, 5, 0) op_6528 (v5842[23:0], v5843[22:0], v6528[27:0]); // 6.0
    wire [21:0] v6529; shift_adder #(20, 20, 1, 1, 22, 1, 0) op_6529 (v5845[19:0], v5846[19:0], v6529[21:0]); // 6.0
    wire [26:0] v6530; shift_adder #(22, 26, 1, 1, 27, -3, 0) op_6530 (v5847[21:0], v5848[25:0], v6530[26:0]); // 6.0
    wire [36:0] v6531; shift_adder #(34, 32, 1, 1, 37, 5, 0) op_6531 (v5849[33:0], v5850[31:0], v6531[36:0]); // 6.0
    wire [33:0] v6532; shift_adder #(32, 28, 1, 1, 34, 6, 0) op_6532 (v5851[31:0], v5852[27:0], v6532[33:0]); // 6.0
    wire [30:0] v6533; shift_adder #(20, 30, 1, 1, 31, -9, 0) op_6533 (v5853[19:0], v5854[29:0], v6533[30:0]); // 6.0
    wire [37:0] v6534; shift_adder #(38, 20, 1, 1, 38, 3, 1) op_6534 (v5855[37:0], v5856[19:0], v6534[37:0]); // 6.0
    wire [33:0] v6535; shift_adder #(33, 30, 1, 1, 34, -1, 0) op_6535 (v5857[32:0], v5858[29:0], v6535[33:0]); // 6.0
    wire [25:0] v6536; shift_adder #(24, 24, 1, 1, 26, -2, 0) op_6536 (v5859[23:0], v5860[23:0], v6536[25:0]); // 6.0
    wire [37:0] v6537; shift_adder #(33, 37, 1, 1, 38, -5, 0) op_6537 (v5861[32:0], v5862[36:0], v6537[37:0]); // 6.0
    wire [38:0] v6538; shift_adder #(38, 31, 1, 1, 39, 7, 0) op_6538 (v5863[37:0], v5864[30:0], v6538[38:0]); // 6.0
    wire [33:0] v6539; shift_adder #(33, 32, 1, 1, 34, -1, 0) op_6539 (v5865[32:0], v5866[31:0], v6539[33:0]); // 6.0
    wire [33:0] v6540; shift_adder #(24, 31, 1, 1, 34, -9, 0) op_6540 (v5867[23:0], v5868[30:0], v6540[33:0]); // 6.0
    wire [27:0] v6541; shift_adder #(22, 28, 1, 1, 28, -2, 0) op_6541 (v5869[21:0], v5870[27:0], v6541[27:0]); // 6.0
    wire [33:0] v6542; shift_adder #(31, 34, 1, 1, 34, -1, 0) op_6542 (v5871[30:0], v5872[33:0], v6542[33:0]); // 6.0
    wire [34:0] v6543; shift_adder #(19, 29, 1, 1, 35, 6, 1) op_6543 (v5873[18:0], v4642[28:0], v6543[34:0]); // 6.0
    wire [33:0] v6544; shift_adder #(32, 27, 1, 1, 34, 6, 0) op_6544 (v5874[31:0], v5875[26:0], v6544[33:0]); // 6.0
    wire [36:0] v6545; shift_adder #(33, 36, 1, 1, 37, -2, 0) op_6545 (v5876[32:0], v5877[35:0], v6545[36:0]); // 6.0
    wire [34:0] v6546; shift_adder #(34, 31, 1, 1, 35, 3, 0) op_6546 (v5878[33:0], v5879[30:0], v6546[34:0]); // 6.0
    wire [37:0] v6547; shift_adder #(35, 21, 1, 1, 38, -3, 1) op_6547 (v5880[34:0], v5881[20:0], v6547[37:0]); // 6.0
    wire [40:0] v6548; shift_adder #(36, 41, 1, 1, 41, -3, 0) op_6548 (v5882[35:0], v5883[40:0], v6548[40:0]); // 6.0
    wire [33:0] v6549; shift_adder #(29, 33, 1, 1, 34, -4, 0) op_6549 (v5884[28:0], v5885[32:0], v6549[33:0]); // 6.0
    wire [33:0] v6550; shift_adder #(29, 32, 1, 1, 34, -5, 0) op_6550 (v5886[28:0], v5887[31:0], v6550[33:0]); // 6.0
    wire [26:0] v6551; shift_adder #(18, 25, 1, 1, 27, -8, 0) op_6551 (v5888[17:0], v5889[24:0], v6551[26:0]); // 6.0
    wire [25:0] v6552; shift_adder #(26, 22, 1, 1, 26, 2, 0) op_6552 (v5890[25:0], v5891[21:0], v6552[25:0]); // 6.0
    wire [32:0] v6553; shift_adder #(29, 25, 1, 1, 33, 7, 0) op_6553 (v5892[28:0], v5893[24:0], v6553[32:0]); // 6.0
    wire [26:0] v6554; shift_adder #(25, 20, 1, 1, 27, 7, 0) op_6554 (v5894[24:0], v5895[19:0], v6554[26:0]); // 6.0
    wire [21:0] v6555; shift_adder #(21, 21, 1, 1, 22, -1, 0) op_6555 (v5896[20:0], v5897[20:0], v6555[21:0]); // 6.0
    wire [37:0] v6556; shift_adder #(33, 35, 1, 1, 38, -4, 0) op_6556 (v5898[32:0], v5899[34:0], v6556[37:0]); // 6.0
    wire [33:0] v6557; shift_adder #(33, 23, 1, 1, 34, 6, 0) op_6557 (v5900[32:0], v5901[22:0], v6557[33:0]); // 6.0
    wire [35:0] v6558; shift_adder #(18, 34, 1, 1, 36, 2, 1) op_6558 (v5902[17:0], v4696[33:0], v6558[35:0]); // 6.0
    wire [36:0] v6559; shift_adder #(24, 37, 1, 1, 37, -12, 0) op_6559 (v5903[23:0], v5904[36:0], v6559[36:0]); // 6.0
    wire [32:0] v6560; shift_adder #(33, 27, 1, 1, 33, 4, 0) op_6560 (v5905[32:0], v5906[26:0], v6560[32:0]); // 6.0
    wire [23:0] v6561; shift_adder #(24, 21, 1, 1, 24, 0, 0) op_6561 (v5907[23:0], v5908[20:0], v6561[23:0]); // 6.0
    wire [32:0] v6562; shift_adder #(32, 20, 1, 1, 33, 12, 0) op_6562 (v5909[31:0], v5910[19:0], v6562[32:0]); // 6.0
    wire [33:0] v6563; shift_adder #(31, 34, 1, 1, 34, -2, 0) op_6563 (v5911[30:0], v5912[33:0], v6563[33:0]); // 6.0
    wire [41:0] v6564; shift_adder #(39, 42, 1, 1, 42, -2, 0) op_6564 (v5913[38:0], v5914[41:0], v6564[41:0]); // 6.0
    wire [21:0] v6565; shift_adder #(20, 19, 1, 1, 22, -2, 0) op_6565 (v5915[19:0], v5916[18:0], v6565[21:0]); // 6.0
    wire [24:0] v6566; shift_adder #(23, 22, 1, 1, 25, 2, 0) op_6566 (v5917[22:0], v5918[21:0], v6566[24:0]); // 6.0
    wire [26:0] v6567; shift_adder #(22, 27, 1, 1, 27, -3, 0) op_6567 (v5919[21:0], v5920[26:0], v6567[26:0]); // 6.0
    wire [28:0] v6568; shift_adder #(26, 25, 1, 1, 29, 4, 0) op_6568 (v5921[25:0], v5922[24:0], v6568[28:0]); // 6.0
    wire [34:0] v6569; shift_adder #(25, 34, 1, 1, 35, -7, 0) op_6569 (v5923[24:0], v5924[33:0], v6569[34:0]); // 6.0
    wire [40:0] v6570; shift_adder #(37, 23, 1, 1, 41, -4, 1) op_6570 (v5925[36:0], v5926[22:0], v6570[40:0]); // 6.0
    wire [23:0] v6571; shift_adder #(24, 20, 1, 1, 24, 0, 0) op_6571 (v5927[23:0], v5928[19:0], v6571[23:0]); // 6.0
    wire [35:0] v6572; shift_adder #(27, 35, 1, 1, 36, -7, 0) op_6572 (v5929[26:0], v5930[34:0], v6572[35:0]); // 6.0
    wire [39:0] v6573; shift_adder #(36, 40, 1, 1, 40, -2, 0) op_6573 (v5931[35:0], v5932[39:0], v6573[39:0]); // 6.0
    wire [36:0] v6574; shift_adder #(35, 35, 1, 1, 37, -1, 0) op_6574 (v5933[34:0], v5934[34:0], v6574[36:0]); // 6.0
    wire [33:0] v6575; shift_adder #(34, 30, 1, 1, 34, 2, 0) op_6575 (v5935[33:0], v5936[29:0], v6575[33:0]); // 6.0
    wire [29:0] v6576; shift_adder #(29, 25, 1, 1, 30, 2, 0) op_6576 (v5937[28:0], v5938[24:0], v6576[29:0]); // 6.0
    wire [27:0] v6577; shift_adder #(27, 26, 1, 1, 28, -1, 0) op_6577 (v5939[26:0], v5940[25:0], v6577[27:0]); // 6.0
    wire [26:0] v6578; shift_adder #(25, 25, 1, 1, 27, 2, 0) op_6578 (v5941[24:0], v5942[24:0], v6578[26:0]); // 6.0
    wire [31:0] v6579; shift_adder #(29, 23, 1, 1, 32, 9, 0) op_6579 (v5943[28:0], v5944[22:0], v6579[31:0]); // 6.0
    wire [34:0] v6580; shift_adder #(33, 35, 1, 1, 35, -1, 0) op_6580 (v5945[32:0], v5946[34:0], v6580[34:0]); // 6.0
    wire [38:0] v6581; shift_adder #(34, 39, 1, 1, 39, -4, 0) op_6581 (v5947[33:0], v5948[38:0], v6581[38:0]); // 6.0
    wire [37:0] v6582; shift_adder #(20, 20, 1, 1, 38, 18, 1) op_6582 (v5949[19:0], v4784[19:0], v6582[37:0]); // 6.0
    wire [36:0] v6583; shift_adder #(31, 19, 1, 1, 37, -6, 1) op_6583 (v5950[30:0], v5951[18:0], v6583[36:0]); // 6.0
    wire [28:0] v6584; shift_adder #(22, 28, 1, 1, 29, -7, 0) op_6584 (v5952[21:0], v5953[27:0], v6584[28:0]); // 6.0
    wire [24:0] v6585; shift_adder #(25, 18, 1, 1, 25, 4, 0) op_6585 (v5954[24:0], v5955[17:0], v6585[24:0]); // 6.0
    wire [27:0] v6586; shift_adder #(25, 27, 1, 1, 28, -2, 0) op_6586 (v5956[24:0], v5957[26:0], v6586[27:0]); // 6.0
    wire [31:0] v6587; shift_adder #(29, 30, 1, 1, 32, -2, 0) op_6587 (v5958[28:0], v5959[29:0], v6587[31:0]); // 6.0
    wire [30:0] v6588; shift_adder #(27, 29, 1, 1, 31, -4, 0) op_6588 (v5960[26:0], v5961[28:0], v6588[30:0]); // 6.0
    wire [30:0] v6589; shift_adder #(26, 29, 1, 1, 31, -4, 0) op_6589 (v5962[25:0], v5963[28:0], v6589[30:0]); // 6.0
    wire [27:0] v6590; shift_adder #(23, 28, 1, 1, 28, -2, 0) op_6590 (v5964[22:0], v5965[27:0], v6590[27:0]); // 6.0
    wire [29:0] v6591; shift_adder #(26, 29, 1, 1, 30, -3, 0) op_6591 (v5773[25:0], v5966[28:0], v6591[29:0]); // 6.0
    wire [27:0] v6592; shift_adder #(26, 26, 1, 1, 28, -2, 0) op_6592 (v5967[25:0], v5968[25:0], v6592[27:0]); // 6.0
    wire [28:0] v6593; shift_adder #(24, 26, 1, 1, 29, -5, 0) op_6593 (v5969[23:0], v5970[25:0], v6593[28:0]); // 6.0
    wire [24:0] v6594; shift_adder #(23, 22, 1, 1, 25, -2, 0) op_6594 (v5971[22:0], v5972[21:0], v6594[24:0]); // 6.0
    wire [26:0] v6595; shift_adder #(25, 23, 1, 1, 27, 4, 0) op_6595 (v5973[24:0], v5974[22:0], v6595[26:0]); // 6.0
    wire [30:0] v6596; shift_adder #(30, 24, 1, 1, 31, 5, 0) op_6596 (v5976[29:0], v5977[23:0], v6596[30:0]); // 6.0
    wire [38:0] v6597; shift_adder #(21, 18, 1, 1, 39, 21, 1) op_6597 (v5978[20:0], v4839[17:0], v6597[38:0]); // 6.0
    wire [30:0] v6598; shift_adder #(24, 30, 1, 1, 31, -5, 0) op_6598 (v5979[23:0], v5980[29:0], v6598[30:0]); // 6.0
    wire [37:0] v6599; shift_adder #(20, 37, 1, 1, 38, -16, 0) op_6599 (v5853[19:0], v5981[36:0], v6599[37:0]); // 6.0
    wire [40:0] v6600; shift_adder #(32, 40, 1, 1, 41, -7, 0) op_6600 (v5982[31:0], v5983[39:0], v6600[40:0]); // 6.0
    wire [40:0] v6601; shift_adder #(41, 19, 1, 1, 41, 1, 1) op_6601 (v5984[40:0], v5985[18:0], v6601[40:0]); // 6.0
    wire [21:0] v6602; shift_adder #(20, 21, 1, 1, 22, 1, 0) op_6602 (v5986[19:0], v5987[20:0], v6602[21:0]); // 6.0
    wire [30:0] v6603; shift_adder #(26, 30, 1, 1, 31, 0, 0) op_6603 (v5988[25:0], v5989[29:0], v6603[30:0]); // 6.0
    wire [27:0] v6604; shift_adder #(25, 24, 1, 1, 28, 4, 0) op_6604 (v5990[24:0], v5991[23:0], v6604[27:0]); // 6.0
    wire [26:0] v6605; shift_adder #(24, 26, 1, 1, 27, -1, 0) op_6605 (v5992[23:0], v5993[25:0], v6605[26:0]); // 6.0
    wire [30:0] v6606; shift_adder #(16, 18, 1, 1, 31, 13, 1) op_6606 (v970[15:0], v5994[17:0], v6606[30:0]); // 6.0
    wire [35:0] v6607; shift_adder #(35, 27, 1, 1, 36, 8, 0) op_6607 (v5995[34:0], v5996[26:0], v6607[35:0]); // 6.0
    wire [38:0] v6608; shift_adder #(20, 27, 1, 1, 39, 12, 1) op_6608 (v5997[19:0], v4876[26:0], v6608[38:0]); // 6.0
    wire [40:0] v6609; shift_adder #(39, 32, 1, 1, 41, 9, 0) op_6609 (v5998[38:0], v5999[31:0], v6609[40:0]); // 6.0
    wire [36:0] v6610; shift_adder #(35, 33, 1, 1, 37, -1, 0) op_6610 (v6000[34:0], v6001[32:0], v6610[36:0]); // 6.0
    wire [31:0] v6611; shift_adder #(30, 30, 1, 1, 32, -1, 0) op_6611 (v6002[29:0], v6003[29:0], v6611[31:0]); // 6.0
    wire [32:0] v6612; shift_adder #(33, 26, 1, 1, 33, 3, 0) op_6612 (v6004[32:0], v6005[25:0], v6612[32:0]); // 6.0
    wire [27:0] v6613; shift_adder #(23, 24, 1, 1, 28, -5, 0) op_6613 (v6006[22:0], v6007[23:0], v6613[27:0]); // 6.0
    wire [25:0] v6614; shift_adder #(23, 21, 1, 1, 26, 5, 0) op_6614 (v6008[22:0], v6009[20:0], v6614[25:0]); // 6.0
    wire [26:0] v6615; shift_adder #(23, 26, 1, 1, 27, -1, 0) op_6615 (v6010[22:0], v6011[25:0], v6615[26:0]); // 6.0
    wire [35:0] v6616; shift_adder #(36, 31, 1, 1, 36, 4, 0) op_6616 (v6012[35:0], v6013[30:0], v6616[35:0]); // 6.0
    wire [37:0] v6617; shift_adder #(35, 29, 1, 1, 38, 8, 0) op_6617 (v6014[34:0], v6015[28:0], v6617[37:0]); // 6.0
    wire [37:0] v6618; shift_adder #(31, 37, 1, 1, 38, -5, 0) op_6618 (v6016[30:0], v6017[36:0], v6618[37:0]); // 6.0
    wire [41:0] v6619; shift_adder #(40, 38, 1, 1, 42, 3, 0) op_6619 (v6018[39:0], v6019[37:0], v6619[41:0]); // 6.0
    wire [23:0] v6620; shift_adder #(24, 20, 1, 1, 24, 0, 0) op_6620 (v6020[23:0], v6021[19:0], v6620[23:0]); // 6.0
    wire [34:0] v6621; shift_adder #(34, 32, 1, 1, 35, 0, 0) op_6621 (v6022[33:0], v6023[31:0], v6621[34:0]); // 6.0
    wire [32:0] v6622; shift_adder #(32, 27, 1, 1, 33, 4, 0) op_6622 (v6024[31:0], v6025[26:0], v6622[32:0]); // 6.0
    wire [31:0] v6623; shift_adder #(27, 31, 1, 1, 32, -4, 0) op_6623 (v6026[26:0], v6027[30:0], v6623[31:0]); // 6.0
    wire [25:0] v6624; shift_adder #(24, 23, 1, 1, 26, -1, 0) op_6624 (v6028[23:0], v6029[22:0], v6624[25:0]); // 6.0
    wire [28:0] v6625; shift_adder #(8, 29, 1, 1, 29, -14, 0) op_6625 (v93[7:0], v6030[28:0], v6625[28:0]); // 6.0
    wire [27:0] v6626; shift_adder #(26, 26, 1, 1, 28, 2, 0) op_6626 (v6031[25:0], v6032[25:0], v6626[27:0]); // 6.0
    wire [35:0] v6627; shift_adder #(36, 32, 1, 1, 36, 1, 0) op_6627 (v6033[35:0], v6034[31:0], v6627[35:0]); // 6.0
    wire [34:0] v6628; shift_adder #(30, 32, 1, 1, 35, -4, 0) op_6628 (v6035[29:0], v6036[31:0], v6628[34:0]); // 6.0
    wire [27:0] v6629; shift_adder #(28, 24, 1, 1, 28, 2, 0) op_6629 (v6037[27:0], v6038[23:0], v6629[27:0]); // 6.0
    wire [30:0] v6630; shift_adder #(27, 26, 1, 1, 31, 4, 0) op_6630 (v6039[26:0], v6040[25:0], v6630[30:0]); // 6.0
    wire [30:0] v6631; shift_adder #(29, 31, 1, 1, 31, 0, 0) op_6631 (v6042[28:0], v6043[30:0], v6631[30:0]); // 6.0
    wire [37:0] v6632; shift_adder #(20, 36, 1, 1, 38, 2, 1) op_6632 (v6044[19:0], v4963[35:0], v6632[37:0]); // 6.0
    wire [35:0] v6633; shift_adder #(32, 35, 1, 1, 36, -2, 0) op_6633 (v6045[31:0], v6046[34:0], v6633[35:0]); // 6.0
    wire [40:0] v6634; shift_adder #(39, 36, 1, 1, 41, 4, 0) op_6634 (v6047[38:0], v6048[35:0], v6634[40:0]); // 6.0
    wire [39:0] v6635; shift_adder #(40, 21, 1, 1, 40, 1, 1) op_6635 (v6049[39:0], v6050[20:0], v6635[39:0]); // 6.0
    wire [27:0] v6636; shift_adder #(23, 26, 1, 1, 28, -4, 0) op_6636 (v6051[22:0], v6052[25:0], v6636[27:0]); // 6.0
    wire [25:0] v6637; shift_adder #(20, 26, 1, 1, 26, -3, 0) op_6637 (v6053[19:0], v6054[25:0], v6637[25:0]); // 6.0
    wire [31:0] v6638; shift_adder #(30, 31, 1, 1, 32, 0, 0) op_6638 (v6055[29:0], v6056[30:0], v6638[31:0]); // 6.0
    wire [31:0] v6639; shift_adder #(31, 28, 1, 1, 32, 3, 0) op_6639 (v6057[30:0], v6058[27:0], v6639[31:0]); // 6.0
    wire [36:0] v6640; shift_adder #(29, 37, 1, 1, 37, -7, 0) op_6640 (v6059[28:0], v6060[36:0], v6640[36:0]); // 6.0
    wire [39:0] v6641; shift_adder #(21, 34, 1, 1, 40, 6, 1) op_6641 (v6061[20:0], v4994[33:0], v6641[39:0]); // 6.0
    wire [39:0] v6642; shift_adder #(31, 39, 1, 1, 40, -9, 0) op_6642 (v6062[30:0], v6063[38:0], v6642[39:0]); // 6.0
    wire [25:0] v6643; shift_adder #(26, 23, 1, 1, 26, 1, 0) op_6643 (v6064[25:0], v6065[22:0], v6643[25:0]); // 6.0
    wire [22:0] v6644; shift_adder #(21, 20, 1, 1, 23, -1, 0) op_6644 (v6066[20:0], v6067[19:0], v6644[22:0]); // 6.0
    wire [28:0] v6645; shift_adder #(28, 27, 1, 1, 29, -1, 0) op_6645 (v6068[27:0], v6069[26:0], v6645[28:0]); // 6.0
    wire [32:0] v6646; shift_adder #(26, 32, 1, 1, 33, -7, 0) op_6646 (v6070[25:0], v6071[31:0], v6646[32:0]); // 6.0
    wire [32:0] v6647; shift_adder #(32, 30, 1, 1, 33, 0, 0) op_6647 (v6072[31:0], v6073[29:0], v6647[32:0]); // 6.0
    wire [27:0] v6648; shift_adder #(27, 27, 1, 1, 28, -1, 0) op_6648 (v6074[26:0], v6075[26:0], v6648[27:0]); // 6.0
    wire [26:0] v6649; shift_adder #(22, 27, 1, 1, 27, -3, 0) op_6649 (v6076[21:0], v6077[26:0], v6649[26:0]); // 6.0
    wire [24:0] v6650; shift_adder #(23, 23, 1, 1, 25, 2, 0) op_6650 (v6078[22:0], v6079[22:0], v6650[24:0]); // 6.0
    wire [31:0] v6651; shift_adder #(30, 28, 1, 1, 32, 3, 0) op_6651 (v6080[29:0], v6081[27:0], v6651[31:0]); // 6.0
    wire [36:0] v6652; shift_adder #(34, 29, 1, 1, 37, 8, 0) op_6652 (v6082[33:0], v6083[28:0], v6652[36:0]); // 6.0
    wire [41:0] v6653; shift_adder #(41, 34, 1, 1, 42, 8, 0) op_6653 (v6084[40:0], v6085[33:0], v6653[41:0]); // 6.0
    wire [27:0] v6654; shift_adder #(28, 22, 1, 1, 28, 4, 0) op_6654 (v6086[27:0], v6087[21:0], v6654[27:0]); // 6.0
    wire [38:0] v6655; shift_adder #(21, 20, 1, 1, 39, 19, 1) op_6655 (v6088[20:0], v5042[19:0], v6655[38:0]); // 6.0
    wire [38:0] v6656; shift_adder #(38, 19, 1, 1, 39, -1, 1) op_6656 (v6089[37:0], v6090[18:0], v6656[38:0]); // 6.0
    wire [35:0] v6657; shift_adder #(35, 25, 1, 1, 36, 9, 0) op_6657 (v6091[34:0], v6092[24:0], v6657[35:0]); // 6.0
    wire [34:0] v6658; shift_adder #(34, 30, 1, 1, 35, 3, 0) op_6658 (v6093[33:0], v6094[29:0], v6658[34:0]); // 6.0
    wire [32:0] v6659; shift_adder #(30, 31, 1, 1, 33, -2, 0) op_6659 (v6095[29:0], v6096[30:0], v6659[32:0]); // 6.0
    wire [26:0] v6660; shift_adder #(27, 23, 1, 1, 27, 1, 0) op_6660 (v6097[26:0], v6098[22:0], v6660[26:0]); // 6.0
    wire [27:0] v6661; shift_adder #(26, 23, 1, 1, 28, 5, 0) op_6661 (v6099[25:0], v6100[22:0], v6661[27:0]); // 6.0
    wire [27:0] v6662; shift_adder #(24, 28, 1, 1, 28, 0, 0) op_6662 (v6101[23:0], v6102[27:0], v6662[27:0]); // 6.0
    wire [33:0] v6663; shift_adder #(33, 27, 1, 1, 34, 6, 0) op_6663 (v6103[32:0], v6104[26:0], v6663[33:0]); // 6.0
    wire [33:0] v6664; shift_adder #(20, 34, 1, 1, 34, -11, 0) op_6664 (v5910[19:0], v6105[33:0], v6664[33:0]); // 6.0
    wire [41:0] v6665; shift_adder #(40, 41, 1, 1, 42, 0, 0) op_6665 (v6106[39:0], v6107[40:0], v6665[41:0]); // 6.0
    wire [26:0] v6666; shift_adder #(26, 22, 1, 1, 27, -1, 0) op_6666 (v6108[25:0], v6109[21:0], v6666[26:0]); // 6.0
    wire [37:0] v6667; shift_adder #(19, 36, 1, 1, 38, 2, 1) op_6667 (v6110[18:0], v5083[35:0], v6667[37:0]); // 6.0
    wire [36:0] v6668; shift_adder #(37, 19, 1, 1, 37, 0, 1) op_6668 (v6111[36:0], v6112[18:0], v6668[36:0]); // 6.0
    wire [35:0] v6669; shift_adder #(34, 34, 1, 1, 36, -1, 0) op_6669 (v6113[33:0], v6114[33:0], v6669[35:0]); // 6.0
    wire [34:0] v6670; shift_adder #(31, 33, 1, 1, 35, -4, 0) op_6670 (v6115[30:0], v6116[32:0], v6670[34:0]); // 6.0
    wire [31:0] v6671; shift_adder #(27, 31, 1, 1, 32, -3, 0) op_6671 (v6117[26:0], v6118[30:0], v6671[31:0]); // 6.0
    wire [30:0] v6672; shift_adder #(24, 29, 1, 1, 31, -7, 0) op_6672 (v6119[23:0], v6120[28:0], v6672[30:0]); // 6.0
    wire [31:0] v6673; shift_adder #(31, 30, 1, 1, 32, 0, 0) op_6673 (v6121[30:0], v6122[29:0], v6673[31:0]); // 6.0
    wire [29:0] v6674; shift_adder #(27, 27, 1, 1, 30, 2, 0) op_6674 (v6123[26:0], v6124[26:0], v6674[29:0]); // 6.0
    wire [26:0] v6675; shift_adder #(23, 27, 1, 1, 27, 0, 0) op_6675 (v6125[22:0], v6126[26:0], v6675[26:0]); // 6.0
    wire [35:0] v6676; shift_adder #(21, 18, 1, 1, 36, 18, 1) op_6676 (v6128[20:0], v5117[17:0], v6676[35:0]); // 6.0
    wire [37:0] v6677; shift_adder #(37, 35, 1, 1, 38, 2, 0) op_6677 (v6129[36:0], v6130[34:0], v6677[37:0]); // 6.0
    wire [42:0] v6678; shift_adder #(38, 42, 1, 1, 43, -2, 0) op_6678 (v6131[37:0], v6132[41:0], v6678[42:0]); // 6.0
    wire [20:0] v6679; shift_adder #(21, 19, 1, 1, 21, 0, 0) op_6679 (v6133[20:0], v6134[18:0], v6679[20:0]); // 6.0
    wire [30:0] v6680; shift_adder #(26, 30, 1, 1, 31, -4, 0) op_6680 (v6135[25:0], v6136[29:0], v6680[30:0]); // 6.0
    wire [29:0] v6681; shift_adder #(30, 27, 1, 1, 30, 1, 0) op_6681 (v6137[29:0], v6138[26:0], v6681[29:0]); // 6.0
    wire [28:0] v6682; shift_adder #(27, 27, 1, 1, 29, -2, 0) op_6682 (v6139[26:0], v6140[26:0], v6682[28:0]); // 6.0
    wire [26:0] v6683; shift_adder #(25, 24, 1, 1, 27, -2, 0) op_6683 (v6141[24:0], v6142[23:0], v6683[26:0]); // 6.0
    wire [23:0] v6684; shift_adder #(22, 23, 1, 1, 24, -1, 0) op_6684 (v6143[21:0], v6144[22:0], v6684[23:0]); // 6.0
    wire [31:0] v6685; shift_adder #(26, 32, 1, 1, 32, -4, 0) op_6685 (v6145[25:0], v6146[31:0], v6685[31:0]); // 6.0
    wire [37:0] v6686; shift_adder #(22, 36, 1, 1, 38, -15, 0) op_6686 (v6147[21:0], v6148[35:0], v6686[37:0]); // 6.0
    wire [32:0] v6687; shift_adder #(27, 32, 1, 1, 33, -6, 0) op_6687 (v6149[26:0], v6150[31:0], v6687[32:0]); // 6.0
    wire [38:0] v6688; shift_adder #(36, 19, 1, 1, 39, -3, 1) op_6688 (v6151[35:0], v6152[18:0], v6688[38:0]); // 6.0
    wire [22:0] v6689; shift_adder #(20, 20, 1, 1, 23, -2, 0) op_6689 (v6153[19:0], v6154[19:0], v6689[22:0]); // 6.0
    wire [30:0] v6690; shift_adder #(27, 29, 1, 1, 31, -3, 0) op_6690 (v6155[26:0], v6156[28:0], v6690[30:0]); // 6.0
    wire [29:0] v6691; shift_adder #(23, 29, 1, 1, 30, -6, 0) op_6691 (v6157[22:0], v6158[28:0], v6691[29:0]); // 6.0
    wire [32:0] v6692; shift_adder #(31, 33, 1, 1, 33, 0, 0) op_6692 (v6159[30:0], v6160[32:0], v6692[32:0]); // 6.0
    wire [33:0] v6693; shift_adder #(32, 33, 1, 1, 34, 0, 0) op_6693 (v5828[31:0], v6161[32:0], v6693[33:0]); // 6.0
    wire [36:0] v6694; shift_adder #(21, 15, 1, 1, 37, 22, 1) op_6694 (v6162[20:0], v5182[14:0], v6694[36:0]); // 6.0
    wire [35:0] v6695; shift_adder #(36, 34, 1, 1, 36, 1, 0) op_6695 (v6163[35:0], v6164[33:0], v6695[35:0]); // 6.0
    wire [29:0] v6696; shift_adder #(26, 26, 1, 1, 30, 4, 0) op_6696 (v6165[25:0], v6166[25:0], v6696[29:0]); // 6.0
    wire [28:0] v6697; shift_adder #(27, 29, 1, 1, 29, -1, 0) op_6697 (v6167[26:0], v6168[28:0], v6697[28:0]); // 6.0
    wire [28:0] v6698; shift_adder #(28, 24, 1, 1, 29, 4, 0) op_6698 (v6169[27:0], v6170[23:0], v6698[28:0]); // 6.0
    wire [34:0] v6699; shift_adder #(35, 28, 1, 1, 35, 5, 0) op_6699 (v6171[34:0], v6172[27:0], v6699[34:0]); // 6.0
    wire [32:0] v6700; shift_adder #(11, 33, 1, 1, 33, -11, 0) op_6700 (v345[10:0], v6173[32:0], v6700[32:0]); // 6.0
    wire [21:0] v6701; shift_adder #(20, 21, 1, 1, 22, 1, 0) op_6701 (v6174[19:0], v6175[20:0], v6701[21:0]); // 6.0
    wire [28:0] v6702; shift_adder #(29, 20, 1, 1, 29, 8, 0) op_6702 (v6177[28:0], v6178[19:0], v6702[28:0]); // 6.0
    wire [28:0] v6703; shift_adder #(26, 26, 1, 1, 29, -3, 0) op_6703 (v6179[25:0], v6180[25:0], v6703[28:0]); // 6.0
    wire [38:0] v6704; shift_adder #(26, 39, 1, 1, 39, -11, 0) op_6704 (v6181[25:0], v6182[38:0], v6704[38:0]); // 6.0
    wire [35:0] v6705; shift_adder #(26, 36, 1, 1, 36, -9, 0) op_6705 (v6183[25:0], v6184[35:0], v6705[35:0]); // 6.0
    wire [38:0] v6706; shift_adder #(39, 19, 1, 1, 39, 2, 1) op_6706 (v6185[38:0], v6186[18:0], v6706[38:0]); // 6.0
    wire [24:0] v6707; shift_adder #(22, 22, 1, 1, 25, -2, 0) op_6707 (v6187[21:0], v6188[21:0], v6707[24:0]); // 6.0
    wire [26:0] v6708; shift_adder #(24, 25, 1, 1, 27, 2, 0) op_6708 (v6189[23:0], v6190[24:0], v6708[26:0]); // 6.0
    wire [29:0] v6709; shift_adder #(27, 27, 1, 1, 30, 3, 0) op_6709 (v6191[26:0], v6192[26:0], v6709[29:0]); // 6.0
    wire [32:0] v6710; shift_adder #(31, 26, 1, 1, 33, 7, 0) op_6710 (v6193[30:0], v5962[25:0], v6710[32:0]); // 6.0
    wire [30:0] v6711; shift_adder #(29, 31, 1, 1, 31, 0, 0) op_6711 (v6194[28:0], v6195[30:0], v6711[30:0]); // 6.0
    wire [36:0] v6712; shift_adder #(19, 21, 1, 1, 37, 16, 1) op_6712 (v6196[18:0], v5243[20:0], v6712[36:0]); // 6.0
    wire [25:0] v6713; shift_adder #(24, 21, 1, 1, 26, -2, 0) op_6713 (v6197[23:0], v6198[20:0], v6713[25:0]); // 6.0
    wire [36:0] v6714; shift_adder #(33, 36, 1, 1, 37, -3, 0) op_6714 (v6199[32:0], v6200[35:0], v6714[36:0]); // 6.0
    wire [38:0] v6715; shift_adder #(37, 39, 1, 1, 39, -1, 0) op_6715 (v6201[36:0], v6202[38:0], v6715[38:0]); // 6.0
    wire [30:0] v6716; shift_adder #(30, 28, 1, 1, 31, 1, 0) op_6716 (v6203[29:0], v6204[27:0], v6716[30:0]); // 6.0
    wire [31:0] v6717; shift_adder #(28, 30, 1, 1, 32, -3, 0) op_6717 (v6205[27:0], v6206[29:0], v6717[31:0]); // 6.0
    wire [30:0] v6718; shift_adder #(31, 26, 1, 1, 31, 3, 0) op_6718 (v6207[30:0], v6208[25:0], v6718[30:0]); // 6.0
    wire [28:0] v6719; shift_adder #(25, 27, 1, 1, 29, -3, 0) op_6719 (v6209[24:0], v6210[26:0], v6719[28:0]); // 6.0
    wire [26:0] v6720; shift_adder #(26, 21, 1, 1, 27, 6, 0) op_6720 (v6211[25:0], v6212[20:0], v6720[26:0]); // 6.0
    wire [26:0] v6721; shift_adder #(25, 26, 1, 1, 27, 1, 0) op_6721 (v6213[24:0], v6214[25:0], v6721[26:0]); // 6.0
    wire [30:0] v6722; shift_adder #(28, 28, 1, 1, 31, 2, 0) op_6722 (v6215[27:0], v6216[27:0], v6722[30:0]); // 6.0
    wire [33:0] v6723; shift_adder #(33, 31, 1, 1, 34, 3, 0) op_6723 (v6217[32:0], v6218[30:0], v6723[33:0]); // 6.0
    wire [40:0] v6724; shift_adder #(37, 40, 1, 1, 41, -2, 0) op_6724 (v6219[36:0], v6220[39:0], v6724[40:0]); // 6.0
    wire [24:0] v6725; shift_adder #(25, 19, 1, 1, 25, 0, 0) op_6725 (v6221[24:0], v6222[18:0], v6725[24:0]); // 6.0
    wire [38:0] v6726; shift_adder #(21, 27, 1, 1, 39, 12, 1) op_6726 (v6223[20:0], v5294[26:0], v6726[38:0]); // 6.0
    wire [34:0] v6727; shift_adder #(34, 28, 1, 1, 35, 6, 0) op_6727 (v6224[33:0], v6225[27:0], v6727[34:0]); // 6.0
    wire [33:0] v6728; shift_adder #(29, 33, 1, 1, 34, -5, 0) op_6728 (v6226[28:0], v6227[32:0], v6728[33:0]); // 6.0
    wire [36:0] v6729; shift_adder #(35, 35, 1, 1, 37, -2, 0) op_6729 (v6228[34:0], v6229[34:0], v6729[36:0]); // 6.0
    wire [29:0] v6730; shift_adder #(25, 28, 1, 1, 30, -4, 0) op_6730 (v6230[24:0], v6231[27:0], v6730[29:0]); // 6.0
    wire [32:0] v6731; shift_adder #(31, 25, 1, 1, 33, 8, 0) op_6731 (v6232[30:0], v6233[24:0], v6731[32:0]); // 6.0
    wire [36:0] v6732; shift_adder #(28, 37, 1, 1, 37, -6, 0) op_6732 (v6234[27:0], v6235[36:0], v6732[36:0]); // 6.0
    wire [26:0] v6733; shift_adder #(20, 27, 1, 1, 27, -2, 0) op_6733 (v6236[19:0], v6237[26:0], v6733[26:0]); // 6.0
    wire [34:0] v6734; shift_adder #(34, 34, 1, 1, 35, 1, 0) op_6734 (v5912[33:0], v6239[33:0], v6734[34:0]); // 6.0
    wire [34:0] v6735; shift_adder #(33, 29, 1, 1, 35, 5, 0) op_6735 (v6240[32:0], v6241[28:0], v6735[34:0]); // 6.0
    wire [40:0] v6736; shift_adder #(40, 39, 1, 1, 41, 2, 0) op_6736 (v6242[39:0], v6243[38:0], v6736[40:0]); // 6.0
    wire [24:0] v6737; shift_adder #(22, 21, 1, 1, 25, -3, 0) op_6737 (v6244[21:0], v6245[20:0], v6737[24:0]); // 6.0
    wire [35:0] v6738; shift_adder #(29, 36, 1, 1, 36, -6, 0) op_6738 (v6042[28:0], v6246[35:0], v6738[35:0]); // 6.0
    wire [33:0] v6739; shift_adder #(33, 29, 1, 1, 34, 2, 0) op_6739 (v6247[32:0], v6248[28:0], v6739[33:0]); // 6.0
    wire [24:0] v6740; shift_adder #(23, 22, 1, 1, 25, -2, 0) op_6740 (v6249[22:0], v6250[21:0], v6740[24:0]); // 6.0
    wire [24:0] v6741; shift_adder #(23, 24, 1, 1, 25, -1, 0) op_6741 (v6251[22:0], v6252[23:0], v6741[24:0]); // 6.0
    wire [25:0] v6742; shift_adder #(22, 21, 1, 1, 26, 5, 0) op_6742 (v6253[21:0], v6254[20:0], v6742[25:0]); // 6.0
    wire [31:0] v6743; shift_adder #(30, 29, 1, 1, 32, 3, 0) op_6743 (v6255[29:0], v6256[28:0], v6743[31:0]); // 6.0
    wire [27:0] v6744; shift_adder #(23, 27, 1, 1, 28, -3, 0) op_6744 (v6257[22:0], v5939[26:0], v6744[27:0]); // 6.0
    wire [32:0] v6745; shift_adder #(27, 32, 1, 1, 33, -4, 0) op_6745 (v6258[26:0], v6259[31:0], v6745[32:0]); // 6.0
    wire [38:0] v6746; shift_adder #(19, 36, 1, 1, 39, 3, 1) op_6746 (v6260[18:0], v5361[35:0], v6746[38:0]); // 6.0
    wire [40:0] v6747; shift_adder #(40, 37, 1, 1, 41, 3, 0) op_6747 (v6261[39:0], v6262[36:0], v6747[40:0]); // 6.0
    wire [26:0] v6748; shift_adder #(27, 22, 1, 1, 27, 3, 0) op_6748 (v6263[26:0], v6264[21:0], v6748[26:0]); // 6.0
    wire [22:0] v6749; shift_adder #(23, 20, 1, 1, 23, 0, 0) op_6749 (v6265[22:0], v6266[19:0], v6749[22:0]); // 6.0
    wire [31:0] v6750; shift_adder #(31, 25, 1, 1, 32, 6, 0) op_6750 (v6267[30:0], v6268[24:0], v6750[31:0]); // 6.0
    wire [30:0] v6751; shift_adder #(19, 30, 1, 1, 31, -11, 0) op_6751 (v6269[18:0], v6270[29:0], v6751[30:0]); // 6.0
    wire [32:0] v6752; shift_adder #(32, 30, 1, 1, 33, 2, 0) op_6752 (v5792[31:0], v6271[29:0], v6752[32:0]); // 6.0
    wire [28:0] v6753; shift_adder #(29, 25, 1, 1, 29, 1, 0) op_6753 (v6272[28:0], v6273[24:0], v6753[28:0]); // 6.0
    wire [26:0] v6754; shift_adder #(23, 27, 1, 1, 27, -1, 0) op_6754 (v6274[22:0], v6275[26:0], v6754[26:0]); // 6.0
    wire [27:0] v6755; shift_adder #(25, 26, 1, 1, 28, 2, 0) op_6755 (v6276[24:0], v6277[25:0], v6755[27:0]); // 6.0
    wire [30:0] v6756; shift_adder #(29, 29, 1, 1, 31, 2, 0) op_6756 (v6278[28:0], v6279[28:0], v6756[30:0]); // 6.0
    wire [37:0] v6757; shift_adder #(33, 38, 1, 1, 38, -2, 0) op_6757 (v6280[32:0], v6281[37:0], v6757[37:0]); // 6.0
    wire [38:0] v6758; shift_adder #(20, 15, 1, 1, 39, 24, 1) op_6758 (v6282[19:0], v5402[14:0], v6758[38:0]); // 6.0
    wire [38:0] v6759; shift_adder #(37, 38, 1, 1, 39, -1, 0) op_6759 (v6283[36:0], v6284[37:0], v6759[38:0]); // 6.0
    wire [24:0] v6760; shift_adder #(22, 23, 1, 1, 25, -3, 0) op_6760 (v6285[21:0], v6286[22:0], v6760[24:0]); // 6.0
    wire [22:0] v6761; shift_adder #(23, 19, 1, 1, 23, 1, 0) op_6761 (v6287[22:0], v6288[18:0], v6761[22:0]); // 6.0
    wire [36:0] v6762; shift_adder #(36, 20, 1, 1, 37, 16, 0) op_6762 (v6289[35:0], v6290[19:0], v6762[36:0]); // 6.0
    wire [34:0] v6763; shift_adder #(35, 30, 1, 1, 35, 3, 0) op_6763 (v6291[34:0], v6292[29:0], v6763[34:0]); // 6.0
    wire [29:0] v6764; shift_adder #(30, 22, 1, 1, 30, 6, 0) op_6764 (v6293[29:0], v6294[21:0], v6764[29:0]); // 6.0
    wire [28:0] v6765; shift_adder #(24, 27, 1, 1, 29, -4, 0) op_6765 (v6295[23:0], v6296[26:0], v6765[28:0]); // 6.0
    wire [27:0] v6766; shift_adder #(25, 28, 1, 1, 28, 0, 0) op_6766 (v6297[24:0], v6298[27:0], v6766[27:0]); // 6.0
    wire [28:0] v6767; shift_adder #(26, 23, 1, 1, 29, 6, 0) op_6767 (v6299[25:0], v6300[22:0], v6767[28:0]); // 6.0
    wire [31:0] v6768; shift_adder #(30, 29, 1, 1, 32, 2, 0) op_6768 (v6301[29:0], v6302[28:0], v6768[31:0]); // 6.0
    wire [34:0] v6769; shift_adder #(34, 32, 1, 1, 35, 3, 0) op_6769 (v6303[33:0], v6304[31:0], v6769[34:0]); // 6.0
    wire [41:0] v6770; shift_adder #(42, 19, 1, 1, 42, 2, 1) op_6770 (v6305[41:0], v6306[18:0], v6770[41:0]); // 6.0
    wire [22:0] v6771; shift_adder #(19, 21, 1, 1, 23, -3, 0) op_6771 (v6307[18:0], v6308[20:0], v6771[22:0]); // 6.0
    wire [36:0] v6772; shift_adder #(20, 28, 1, 1, 37, 9, 1) op_6772 (v6309[19:0], v5450[27:0], v6772[36:0]); // 6.0
    wire [37:0] v6773; shift_adder #(37, 36, 1, 1, 38, 1, 0) op_6773 (v6310[36:0], v6311[35:0], v6773[37:0]); // 6.0
    wire [33:0] v6774; shift_adder #(33, 29, 1, 1, 34, 3, 0) op_6774 (v6312[32:0], v6313[28:0], v6774[33:0]); // 6.0
    wire [31:0] v6775; shift_adder #(31, 24, 1, 1, 32, 7, 0) op_6775 (v6314[30:0], v5977[23:0], v6775[31:0]); // 6.0
    wire [32:0] v6776; shift_adder #(32, 29, 1, 1, 33, -1, 0) op_6776 (v6315[31:0], v6316[28:0], v6776[32:0]); // 6.0
    wire [27:0] v6777; shift_adder #(26, 23, 1, 1, 28, -2, 0) op_6777 (v6317[25:0], v6318[22:0], v6777[27:0]); // 6.0
    wire [23:0] v6778; shift_adder #(19, 24, 1, 1, 24, 0, 0) op_6778 (v6319[18:0], v6320[23:0], v6778[23:0]); // 6.0
    wire [33:0] v6779; shift_adder #(25, 34, 1, 1, 34, -6, 0) op_6779 (v6321[24:0], v6322[33:0], v6779[33:0]); // 6.0
    wire [32:0] v6780; shift_adder #(28, 32, 1, 1, 33, -5, 0) op_6780 (v6323[27:0], v6324[31:0], v6780[32:0]); // 6.0
    wire [34:0] v6781; shift_adder #(25, 35, 1, 1, 35, -8, 0) op_6781 (v6209[24:0], v6325[34:0], v6781[34:0]); // 6.0
    wire [39:0] v6782; shift_adder #(29, 39, 1, 1, 40, -10, 0) op_6782 (v6326[28:0], v6327[38:0], v6782[39:0]); // 6.0
    wire [38:0] v6783; shift_adder #(37, 37, 1, 1, 39, 1, 0) op_6783 (v6328[36:0], v6329[36:0], v6783[38:0]); // 6.0
    wire [21:0] v6784; shift_adder #(22, 19, 1, 1, 22, 0, 0) op_6784 (v6330[21:0], v6331[18:0], v6784[21:0]); // 6.0
    wire [31:0] v6785; shift_adder #(32, 28, 1, 1, 32, 1, 0) op_6785 (v6332[31:0], v6333[27:0], v6785[31:0]); // 6.0
    wire [30:0] v6786; shift_adder #(29, 29, 1, 1, 31, -2, 0) op_6786 (v6334[28:0], v6335[28:0], v6786[30:0]); // 6.0
    wire [29:0] v6787; shift_adder #(22, 28, 1, 1, 30, -8, 0) op_6787 (v6143[21:0], v6336[27:0], v6787[29:0]); // 6.0
    wire [25:0] v6788; shift_adder #(25, 22, 1, 1, 26, 1, 0) op_6788 (v6337[24:0], v6338[21:0], v6788[25:0]); // 6.0
    wire [27:0] v6789; shift_adder #(24, 23, 1, 1, 28, 5, 0) op_6789 (v6339[23:0], v6340[22:0], v6789[27:0]); // 6.0
    wire [25:0] v6790; shift_adder #(21, 25, 1, 1, 26, -3, 0) op_6790 (v6341[20:0], v6342[24:0], v6790[25:0]); // 6.0
    wire [32:0] v6791; shift_adder #(27, 33, 1, 1, 33, -4, 0) op_6791 (v6343[26:0], v6344[32:0], v6791[32:0]); // 6.0
    wire [36:0] v6792; shift_adder #(35, 31, 1, 1, 37, 5, 0) op_6792 (v6345[34:0], v6118[30:0], v6792[36:0]); // 6.0
    wire [38:0] v6793; shift_adder #(39, 18, 1, 1, 39, 4, 1) op_6793 (v6346[38:0], v5802[17:0], v6793[38:0]); // 6.0
    wire [25:0] v6794; shift_adder #(26, 23, 1, 1, 26, 1, 0) op_6794 (v6347[25:0], v6348[22:0], v6794[25:0]); // 6.0
    wire [37:0] v6795; shift_adder #(34, 38, 1, 1, 38, -2, 0) op_6795 (v6349[33:0], v6350[37:0], v6795[37:0]); // 6.0
    wire [41:0] v6796; shift_adder #(33, 41, 1, 1, 42, -7, 0) op_6796 (v6351[32:0], v6352[40:0], v6796[41:0]); // 6.0
    wire [32:0] v6797; shift_adder #(33, 29, 1, 1, 33, 3, 0) op_6797 (v6353[32:0], v6354[28:0], v6797[32:0]); // 6.0
    wire [34:0] v6798; shift_adder #(34, 31, 1, 1, 35, 2, 0) op_6798 (v6355[33:0], v6356[30:0], v6798[34:0]); // 6.0
    wire [32:0] v6799; shift_adder #(33, 30, 1, 1, 33, 1, 0) op_6799 (v6357[32:0], v6358[29:0], v6799[32:0]); // 6.0
    wire [28:0] v6800; shift_adder #(29, 24, 1, 1, 29, 1, 0) op_6800 (v6359[28:0], v6360[23:0], v6800[28:0]); // 6.0
    wire [27:0] v6801; shift_adder #(25, 26, 1, 1, 28, 2, 0) op_6801 (v6361[24:0], v6362[25:0], v6801[27:0]); // 6.0
    wire [31:0] v6802; shift_adder #(31, 20, 1, 1, 32, 11, 0) op_6802 (v6363[30:0], v6364[19:0], v6802[31:0]); // 6.0
    wire [29:0] v6803; shift_adder #(29, 28, 1, 1, 30, 0, 0) op_6803 (v6365[28:0], v6366[27:0], v6803[29:0]); // 6.0
    wire [30:0] v6804; shift_adder #(26, 29, 1, 1, 31, -5, 0) op_6804 (v6367[25:0], v6368[28:0], v6804[30:0]); // 6.0
    wire [34:0] v6805; shift_adder #(32, 30, 1, 1, 35, 5, 0) op_6805 (v6369[31:0], v6370[29:0], v6805[34:0]); // 6.0
    wire [35:0] v6806; shift_adder #(34, 36, 1, 1, 36, 0, 0) op_6806 (v6371[33:0], v6372[35:0], v6806[35:0]); // 6.0
    wire [39:0] v6807; shift_adder #(24, 35, 1, 1, 40, 5, 1) op_6807 (v6373[23:0], v5562[34:0], v6807[39:0]); // 6.0
    wire [41:0] v6808; shift_adder #(33, 41, 1, 1, 42, -7, 0) op_6808 (v6374[32:0], v6375[40:0], v6808[41:0]); // 6.0
    wire [39:0] v6809; shift_adder #(40, 18, 1, 1, 40, 2, 1) op_6809 (v6376[39:0], v6377[17:0], v6809[39:0]); // 6.0
    wire [30:0] v6810; shift_adder #(23, 26, 1, 1, 31, -8, 0) op_6810 (v6378[22:0], v6379[25:0], v6810[30:0]); // 6.0
    wire [22:0] v6811; shift_adder #(23, 18, 1, 1, 23, 2, 0) op_6811 (v6380[22:0], v6381[17:0], v6811[22:0]); // 6.0
    wire [23:0] v6812; shift_adder #(21, 23, 1, 1, 24, -1, 0) op_6812 (v6382[20:0], v6383[22:0], v6812[23:0]); // 6.0
    wire [26:0] v6813; shift_adder #(24, 26, 1, 1, 27, 1, 0) op_6813 (v6384[23:0], v6385[25:0], v6813[26:0]); // 6.0
    wire [31:0] v6814; shift_adder #(30, 31, 1, 1, 32, 1, 0) op_6814 (v6386[29:0], v6387[30:0], v6814[31:0]); // 6.0
    wire [31:0] v6815; shift_adder #(29, 32, 1, 1, 32, -2, 0) op_6815 (v6388[28:0], v6389[31:0], v6815[31:0]); // 6.0
    wire [39:0] v6816; shift_adder #(37, 23, 1, 1, 40, 16, 0) op_6816 (v6390[36:0], v6391[22:0], v6816[39:0]); // 6.0
    wire [39:0] v6817; shift_adder #(37, 39, 1, 1, 40, -1, 0) op_6817 (v6392[36:0], v6393[38:0], v6817[39:0]); // 6.0
    wire [38:0] v6818; shift_adder #(39, 21, 1, 1, 39, 1, 1) op_6818 (v6394[38:0], v6395[20:0], v6818[38:0]); // 6.0
    wire [35:0] v6819; shift_adder #(35, 29, 1, 1, 36, 5, 0) op_6819 (v6396[34:0], v6397[28:0], v6819[35:0]); // 6.0
    wire [30:0] v6820; shift_adder #(28, 28, 1, 1, 31, -2, 0) op_6820 (v6398[27:0], v6399[27:0], v6820[30:0]); // 6.0
    wire [28:0] v6821; shift_adder #(23, 27, 1, 1, 29, -5, 0) op_6821 (v6400[22:0], v6401[26:0], v6821[28:0]); // 6.0
    wire [25:0] v6822; shift_adder #(25, 21, 1, 1, 26, 3, 0) op_6822 (v6402[24:0], v6403[20:0], v6822[25:0]); // 6.0
    wire [29:0] v6823; shift_adder #(23, 30, 1, 1, 30, -3, 0) op_6823 (v6404[22:0], v6405[29:0], v6823[29:0]); // 6.0
    wire [33:0] v6824; shift_adder #(33, 25, 1, 1, 34, 9, 0) op_6824 (v6406[32:0], v6407[24:0], v6824[33:0]); // 6.0
    wire [27:0] v6825; shift_adder #(26, 25, 1, 1, 28, 3, 0) op_6825 (v6408[25:0], v6409[24:0], v6825[27:0]); // 6.0
    wire [40:0] v6826; shift_adder #(38, 40, 1, 1, 41, -2, 0) op_6826 (v6411[37:0], v6412[39:0], v6826[40:0]); // 6.0
    wire [23:0] v6827; shift_adder #(20, 22, 1, 1, 24, -4, 0) op_6827 (v6413[19:0], v6414[21:0], v6827[23:0]); // 6.0
    wire [41:0] v6828; shift_adder #(30, 42, 1, 1, 42, -10, 0) op_6828 (v6415[29:0], v6416[41:0], v6828[41:0]); // 6.0
    wire [35:0] v6829; shift_adder #(19, 23, 1, 1, 36, 13, 1) op_6829 (v6417[18:0], v5639[22:0], v6829[35:0]); // 6.0
    wire [35:0] v6830; shift_adder #(33, 33, 1, 1, 36, -2, 0) op_6830 (v6418[32:0], v6419[32:0], v6830[35:0]); // 6.0
    wire [31:0] v6831; shift_adder #(26, 31, 1, 1, 32, -6, 0) op_6831 (v6420[25:0], v6421[30:0], v6831[31:0]); // 6.0
    wire [32:0] v6832; shift_adder #(30, 31, 1, 1, 33, -2, 0) op_6832 (v6422[29:0], v6423[30:0], v6832[32:0]); // 6.0
    wire [28:0] v6833; shift_adder #(28, 22, 1, 1, 29, 6, 0) op_6833 (v6424[27:0], v6425[21:0], v6833[28:0]); // 6.0
    wire [21:0] v6834; shift_adder #(20, 20, 1, 1, 22, 2, 0) op_6834 (v6426[19:0], v6427[19:0], v6834[21:0]); // 6.0
    wire [27:0] v6835; shift_adder #(25, 25, 1, 1, 28, 3, 0) op_6835 (v6428[24:0], v6429[24:0], v6835[27:0]); // 6.0
    wire [33:0] v6836; shift_adder #(32, 33, 1, 1, 34, -2, 0) op_6836 (v6430[31:0], v6431[32:0], v6836[33:0]); // 6.0
    wire [32:0] v6837; shift_adder #(30, 32, 1, 1, 33, 1, 0) op_6837 (v6432[29:0], v6433[31:0], v6837[32:0]); // 6.0
    wire [34:0] v6838; shift_adder #(33, 26, 1, 1, 35, 8, 0) op_6838 (v6434[32:0], v6435[25:0], v6838[34:0]); // 6.0
    wire [32:0] v6839; shift_adder #(33, 31, 1, 1, 33, 1, 0) op_6839 (v6436[32:0], v6437[30:0], v6839[32:0]); // 6.0
    wire [39:0] v6840; shift_adder #(31, 39, 1, 1, 40, -7, 0) op_6840 (v6438[30:0], v6439[38:0], v6840[39:0]); // 6.0
    wire [32:0] v6841; shift_adder #(32, 31, 1, 1, 33, -1, 0) op_6841 (v6440[31:0], v6441[30:0], v6841[32:0]); // 6.0
    wire [31:0] v6842; shift_adder #(26, 30, 1, 1, 32, -6, 0) op_6842 (v6442[25:0], v6443[29:0], v6842[31:0]); // 6.0
    wire [26:0] v6843; shift_adder #(23, 24, 1, 1, 27, -3, 0) op_6843 (v6444[22:0], v6445[23:0], v6843[26:0]); // 6.0
    wire [19:0] v6844; shift_adder #(20, 17, 1, 1, 20, 0, 0) op_6844 (v6446[19:0], v6447[16:0], v6844[19:0]); // 6.0
    wire [23:0] v6845; shift_adder #(21, 23, 1, 1, 24, -2, 0) op_6845 (v6448[20:0], v6449[22:0], v6845[23:0]); // 6.0
    wire [25:0] v6846; shift_adder #(25, 24, 1, 1, 26, 2, 0) op_6846 (v6450[24:0], v6451[23:0], v6846[25:0]); // 6.0
    wire [33:0] v6847; shift_adder #(27, 32, 1, 1, 34, -7, 0) op_6847 (v6452[26:0], v6453[31:0], v6847[33:0]); // 6.0
    wire [31:0] v6848; shift_adder #(27, 31, 1, 1, 32, -2, 0) op_6848 (v6454[26:0], v6455[30:0], v6848[31:0]); // 6.0
    wire [32:0] v6849; shift_adder #(25, 33, 1, 1, 33, -6, 0) op_6849 (v6456[24:0], v6457[32:0], v6849[32:0]); // 6.0
    wire [35:0] v6850; shift_adder #(34, 35, 1, 1, 36, 0, 0) op_6850 (v6458[33:0], v6459[34:0], v6850[35:0]); // 6.0
    wire [41:0] v6851; shift_adder #(41, 39, 1, 1, 42, 3, 0) op_6851 (v6460[40:0], v6461[38:0], v6851[41:0]); // 6.0
    wire [34:0] v6852; shift_adder #(28, 34, 1, 1, 35, -7, 0) op_6852 (v6462[27:0], v6463[33:0], v6852[34:0]); // 6.0
    wire [31:0] v6853; shift_adder #(27, 29, 1, 1, 32, -5, 0) op_6853 (v6464[26:0], v6465[28:0], v6853[31:0]); // 6.0
    wire [28:0] v6854; shift_adder #(29, 26, 1, 1, 29, 0, 0) op_6854 (v6466[28:0], v6467[25:0], v6854[28:0]); // 6.0
    wire [24:0] v6855; shift_adder #(20, 22, 1, 1, 25, -5, 0) op_6855 (v6468[19:0], v6469[21:0], v6855[24:0]); // 6.0
    wire [33:0] v6856; shift_adder #(30, 30, 1, 1, 34, 4, 0) op_6856 (v6470[29:0], v6471[29:0], v6856[33:0]); // 6.0
    wire [30:0] v6857; shift_adder #(27, 29, 1, 1, 31, -3, 0) op_6857 (v6472[26:0], v5961[28:0], v6857[30:0]); // 6.0
    wire [26:0] v6858; shift_adder #(24, 23, 1, 1, 27, 3, 0) op_6858 (v6473[23:0], v6474[22:0], v6858[26:0]); // 6.0
    wire [33:0] v6859; shift_adder #(22, 34, 1, 1, 34, -11, 0) op_6859 (v6264[21:0], v6476[33:0], v6859[33:0]); // 6.0
    wire [38:0] v6860; shift_adder #(39, 21, 1, 1, 39, 0, 1) op_6860 (v6477[38:0], v6478[20:0], v6860[38:0]); // 6.0
    wire [37:0] v6861; shift_adder #(24, 37, 1, 1, 38, -13, 0) op_6861 (v6479[23:0], v6480[36:0], v6861[37:0]); // 6.0
    wire [37:0] v6862; shift_adder #(28, 38, 1, 1, 38, -8, 0) op_6862 (v6481[27:0], v6482[37:0], v6862[37:0]); // 6.0
    wire [38:0] v6863; shift_adder #(34, 39, 1, 1, 39, -3, 0) op_6863 (v6483[33:0], v6484[38:0], v6863[38:0]); // 6.0
    wire [30:0] v6864; shift_adder #(27, 29, 1, 1, 31, -4, 0) op_6864 (v6485[26:0], v6486[28:0], v6864[30:0]); // 6.0
    wire [34:0] v6865; shift_adder #(35, 30, 1, 1, 35, 1, 0) op_6865 (v6487[34:0], v6488[29:0], v6865[34:0]); // 6.0
    wire [26:0] v6866; shift_adder #(25, 24, 1, 1, 27, -2, 0) op_6866 (v6489[24:0], v6490[23:0], v6866[26:0]); // 6.0
    wire [29:0] v6867; shift_adder #(26, 30, 1, 1, 30, 0, 0) op_6867 (v6491[25:0], v6492[29:0], v6867[29:0]); // 7.0
    wire [33:0] v6868; shift_adder #(33, 32, 1, 1, 34, 1, 0) op_6868 (v6493[32:0], v6494[31:0], v6868[33:0]); // 7.0
    wire [34:0] v6869; shift_adder #(30, 33, 1, 1, 35, -5, 0) op_6869 (v6495[29:0], v6496[32:0], v6869[34:0]); // 7.0
    wire [38:0] v6870; shift_adder #(38, 30, 1, 1, 39, 8, 0) op_6870 (v6497[37:0], v6498[29:0], v6870[38:0]); // 7.0
    wire [39:0] v6871; shift_adder #(26, 32, 1, 1, 40, 8, 1) op_6871 (v6499[25:0], v5787[31:0], v6871[39:0]); // 7.0
    wire [37:0] v6872; shift_adder #(38, 23, 1, 1, 38, 0, 1) op_6872 (v6500[37:0], v6501[22:0], v6872[37:0]); // 7.0
    wire [32:0] v6873; shift_adder #(33, 25, 1, 1, 33, 4, 0) op_6873 (v6502[32:0], v6503[24:0], v6873[32:0]); // 7.0
    wire [31:0] v6874; shift_adder #(26, 30, 1, 1, 32, 2, 0) op_6874 (v6504[25:0], v6505[29:0], v6874[31:0]); // 7.0
    wire [32:0] v6875; shift_adder #(24, 30, 1, 1, 33, -8, 0) op_6875 (v6507[23:0], v6508[29:0], v6875[32:0]); // 7.0
    wire [35:0] v6876; shift_adder #(34, 35, 1, 1, 36, 0, 0) op_6876 (v6509[33:0], v6510[34:0], v6876[35:0]); // 7.0
    wire [37:0] v6877; shift_adder #(37, 25, 1, 1, 38, -1, 1) op_6877 (v6511[36:0], v6512[24:0], v6877[37:0]); // 7.0
    wire [40:0] v6878; shift_adder #(38, 41, 1, 1, 41, -2, 0) op_6878 (v6513[37:0], v6514[40:0], v6878[40:0]); // 7.0
    wire [31:0] v6879; shift_adder #(30, 27, 1, 1, 32, -2, 0) op_6879 (v6515[29:0], v6516[26:0], v6879[31:0]); // 7.0
    wire [33:0] v6880; shift_adder #(31, 31, 1, 1, 34, 3, 0) op_6880 (v6517[30:0], v6518[30:0], v6880[33:0]); // 7.0
    wire [33:0] v6881; shift_adder #(25, 33, 1, 1, 34, -8, 0) op_6881 (v6520[24:0], v6521[32:0], v6881[33:0]); // 7.0
    wire [40:0] v6882; shift_adder #(41, 38, 1, 1, 41, 2, 0) op_6882 (v6522[40:0], v6523[37:0], v6882[40:0]); // 7.0
    wire [31:0] v6883; shift_adder #(32, 22, 1, 1, 32, 6, 0) op_6883 (v6524[31:0], v6525[21:0], v6883[31:0]); // 7.0
    wire [35:0] v6884; shift_adder #(33, 35, 1, 1, 36, 1, 0) op_6884 (v6526[32:0], v6527[34:0], v6884[35:0]); // 7.0
    wire [43:0] v6885; shift_adder #(28, 38, 1, 1, 44, 6, 1) op_6885 (v6528[27:0], v5844[37:0], v6885[43:0]); // 7.0
    wire [28:0] v6886; shift_adder #(22, 27, 1, 1, 29, 2, 0) op_6886 (v6529[21:0], v6530[26:0], v6886[28:0]); // 7.0
    wire [39:0] v6887; shift_adder #(37, 34, 1, 1, 40, 6, 0) op_6887 (v6531[36:0], v6532[33:0], v6887[39:0]); // 7.0
    wire [38:0] v6888; shift_adder #(31, 38, 1, 1, 39, -7, 0) op_6888 (v6533[30:0], v6534[37:0], v6888[38:0]); // 7.0
    wire [33:0] v6889; shift_adder #(34, 26, 1, 1, 34, 2, 0) op_6889 (v6535[33:0], v6536[25:0], v6889[33:0]); // 7.0
    wire [39:0] v6890; shift_adder #(38, 39, 1, 1, 40, -1, 0) op_6890 (v6537[37:0], v6538[38:0], v6890[39:0]); // 7.0
    wire [35:0] v6891; shift_adder #(34, 34, 1, 1, 36, -2, 0) op_6891 (v6539[33:0], v6540[33:0], v6891[35:0]); // 7.0
    wire [33:0] v6892; shift_adder #(28, 34, 1, 1, 34, -2, 0) op_6892 (v6541[27:0], v6542[33:0], v6892[33:0]); // 7.0
    wire [35:0] v6893; shift_adder #(35, 34, 1, 1, 36, 1, 0) op_6893 (v6543[34:0], v6544[33:0], v6893[35:0]); // 7.0
    wire [38:0] v6894; shift_adder #(37, 35, 1, 1, 39, 3, 0) op_6894 (v6545[36:0], v6546[34:0], v6894[38:0]); // 7.0
    wire [41:0] v6895; shift_adder #(38, 41, 1, 1, 42, -2, 0) op_6895 (v6547[37:0], v6548[40:0], v6895[41:0]); // 7.0
    wire [36:0] v6896; shift_adder #(34, 34, 1, 1, 37, -2, 0) op_6896 (v6549[33:0], v6550[33:0], v6896[36:0]); // 7.0
    wire [29:0] v6897; shift_adder #(27, 26, 1, 1, 30, -3, 0) op_6897 (v6551[26:0], v6552[25:0], v6897[29:0]); // 7.0
    wire [36:0] v6898; shift_adder #(33, 27, 1, 1, 37, 10, 0) op_6898 (v6553[32:0], v6554[26:0], v6898[36:0]); // 7.0
    wire [37:0] v6899; shift_adder #(38, 34, 1, 1, 38, 2, 0) op_6899 (v6556[37:0], v6557[33:0], v6899[37:0]); // 7.0
    wire [37:0] v6900; shift_adder #(36, 37, 1, 1, 38, 0, 0) op_6900 (v6558[35:0], v6559[36:0], v6900[37:0]); // 7.0
    wire [32:0] v6901; shift_adder #(33, 24, 1, 1, 33, 5, 0) op_6901 (v6560[32:0], v6561[23:0], v6901[32:0]); // 7.0
    wire [36:0] v6902; shift_adder #(33, 34, 1, 1, 37, 2, 0) op_6902 (v6562[32:0], v6563[33:0], v6902[36:0]); // 7.0
    wire [41:0] v6903; shift_adder #(42, 22, 1, 1, 42, 3, 1) op_6903 (v6564[41:0], v6565[21:0], v6903[41:0]); // 7.0
    wire [27:0] v6904; shift_adder #(25, 27, 1, 1, 28, 1, 0) op_6904 (v6566[24:0], v6567[26:0], v6904[27:0]); // 7.0
    wire [34:0] v6905; shift_adder #(29, 35, 1, 1, 35, -2, 0) op_6905 (v6568[28:0], v6569[34:0], v6905[34:0]); // 7.0
    wire [40:0] v6906; shift_adder #(41, 24, 1, 1, 41, 5, 1) op_6906 (v6570[40:0], v6571[23:0], v6906[40:0]); // 7.0
    wire [40:0] v6907; shift_adder #(36, 40, 1, 1, 41, -3, 0) op_6907 (v6572[35:0], v6573[39:0], v6907[40:0]); // 7.0
    wire [36:0] v6908; shift_adder #(37, 34, 1, 1, 37, 0, 0) op_6908 (v6574[36:0], v6575[33:0], v6908[36:0]); // 7.0
    wire [30:0] v6909; shift_adder #(30, 28, 1, 1, 31, -1, 0) op_6909 (v6576[29:0], v6577[27:0], v6909[30:0]); // 7.0
    wire [31:0] v6910; shift_adder #(27, 32, 1, 1, 32, -1, 0) op_6910 (v6578[26:0], v6579[31:0], v6910[31:0]); // 7.0
    wire [39:0] v6911; shift_adder #(35, 39, 1, 1, 40, -3, 0) op_6911 (v6580[34:0], v6581[38:0], v6911[39:0]); // 7.0
    wire [38:0] v6912; shift_adder #(38, 37, 1, 1, 39, 1, 0) op_6912 (v6582[37:0], v6583[36:0], v6912[38:0]); // 7.0
    wire [30:0] v6913; shift_adder #(29, 25, 1, 1, 31, -1, 0) op_6913 (v6584[28:0], v6585[24:0], v6913[30:0]); // 7.0
    wire [33:0] v6914; shift_adder #(28, 32, 1, 1, 34, -6, 0) op_6914 (v6586[27:0], v6587[31:0], v6914[33:0]); // 7.0
    wire [31:0] v6915; shift_adder #(31, 31, 1, 1, 32, 0, 0) op_6915 (v6588[30:0], v6589[30:0], v6915[31:0]); // 7.0
    wire [29:0] v6916; shift_adder #(28, 30, 1, 1, 30, 0, 0) op_6916 (v6590[27:0], v6591[29:0], v6916[29:0]); // 7.0
    wire [30:0] v6917; shift_adder #(29, 25, 1, 1, 31, -2, 0) op_6917 (v6593[28:0], v6594[24:0], v6917[30:0]); // 7.0
    wire [39:0] v6918; shift_adder #(27, 26, 1, 1, 40, 14, 1) op_6918 (v6595[26:0], v5975[25:0], v6918[39:0]); // 7.0
    wire [38:0] v6919; shift_adder #(31, 39, 1, 1, 39, -6, 0) op_6919 (v6596[30:0], v6597[38:0], v6919[38:0]); // 7.0
    wire [38:0] v6920; shift_adder #(31, 38, 1, 1, 39, -7, 0) op_6920 (v6598[30:0], v6599[37:0], v6920[38:0]); // 7.0
    wire [41:0] v6921; shift_adder #(41, 41, 1, 1, 42, 0, 0) op_6921 (v6600[40:0], v6601[40:0], v6921[41:0]); // 7.0
    wire [30:0] v6922; shift_adder #(22, 31, 1, 1, 31, -3, 0) op_6922 (v6602[21:0], v6603[30:0], v6922[30:0]); // 7.0
    wire [29:0] v6923; shift_adder #(28, 27, 1, 1, 30, 3, 0) op_6923 (v6604[27:0], v6605[26:0], v6923[29:0]); // 7.0
    wire [36:0] v6924; shift_adder #(31, 36, 1, 1, 37, -4, 0) op_6924 (v6606[30:0], v6607[35:0], v6924[36:0]); // 7.0
    wire [41:0] v6925; shift_adder #(39, 41, 1, 1, 42, -1, 0) op_6925 (v6608[38:0], v6609[40:0], v6925[41:0]); // 7.0
    wire [36:0] v6926; shift_adder #(37, 32, 1, 1, 37, 1, 0) op_6926 (v6610[36:0], v6611[31:0], v6926[36:0]); // 7.0
    wire [34:0] v6927; shift_adder #(33, 28, 1, 1, 35, -2, 0) op_6927 (v6612[32:0], v6613[27:0], v6927[34:0]); // 7.0
    wire [31:0] v6928; shift_adder #(26, 27, 1, 1, 32, 5, 0) op_6928 (v6614[25:0], v6615[26:0], v6928[31:0]); // 7.0
    wire [39:0] v6929; shift_adder #(38, 38, 1, 1, 40, 2, 0) op_6929 (v6617[37:0], v6618[37:0], v6929[39:0]); // 7.0
    wire [41:0] v6930; shift_adder #(42, 24, 1, 1, 42, 2, 1) op_6930 (v6619[41:0], v6620[23:0], v6930[41:0]); // 7.0
    wire [35:0] v6931; shift_adder #(35, 33, 1, 1, 36, -1, 0) op_6931 (v6621[34:0], v6622[32:0], v6931[35:0]); // 7.0
    wire [31:0] v6932; shift_adder #(32, 26, 1, 1, 32, 3, 0) op_6932 (v6623[31:0], v6624[25:0], v6932[31:0]); // 7.0
    wire [30:0] v6933; shift_adder #(29, 28, 1, 1, 31, 2, 0) op_6933 (v6625[28:0], v6626[27:0], v6933[30:0]); // 7.0
    wire [34:0] v6934; shift_adder #(35, 28, 1, 1, 35, 2, 0) op_6934 (v6628[34:0], v6629[27:0], v6934[34:0]); // 7.0
    wire [37:0] v6935; shift_adder #(31, 34, 1, 1, 38, 4, 1) op_6935 (v6630[30:0], v6041[33:0], v6935[37:0]); // 7.0
    wire [37:0] v6936; shift_adder #(31, 38, 1, 1, 38, -4, 0) op_6936 (v6631[30:0], v6632[37:0], v6936[37:0]); // 7.0
    wire [40:0] v6937; shift_adder #(36, 41, 1, 1, 41, -4, 0) op_6937 (v6633[35:0], v6634[40:0], v6937[40:0]); // 7.0
    wire [40:0] v6938; shift_adder #(40, 28, 1, 1, 41, -1, 1) op_6938 (v6635[39:0], v6636[27:0], v6938[40:0]); // 7.0
    wire [31:0] v6939; shift_adder #(26, 32, 1, 1, 32, -1, 0) op_6939 (v6637[25:0], v6638[31:0], v6939[31:0]); // 7.0
    wire [37:0] v6940; shift_adder #(32, 37, 1, 1, 38, -4, 0) op_6940 (v6639[31:0], v6640[36:0], v6940[37:0]); // 7.0
    wire [41:0] v6941; shift_adder #(40, 40, 1, 1, 42, 1, 0) op_6941 (v6641[39:0], v6642[39:0], v6941[41:0]); // 7.0
    wire [26:0] v6942; shift_adder #(26, 23, 1, 1, 27, -1, 0) op_6942 (v6643[25:0], v6644[22:0], v6942[26:0]); // 7.0
    wire [35:0] v6943; shift_adder #(29, 33, 1, 1, 36, -7, 0) op_6943 (v6645[28:0], v6646[32:0], v6943[35:0]); // 7.0
    wire [32:0] v6944; shift_adder #(33, 28, 1, 1, 33, 0, 0) op_6944 (v6647[32:0], v6648[27:0], v6944[32:0]); // 7.0
    wire [31:0] v6945; shift_adder #(27, 25, 1, 1, 32, 6, 0) op_6945 (v6649[26:0], v6650[24:0], v6945[31:0]); // 7.0
    wire [36:0] v6946; shift_adder #(32, 37, 1, 1, 37, -2, 0) op_6946 (v6651[31:0], v6652[36:0], v6946[36:0]); // 7.0
    wire [42:0] v6947; shift_adder #(42, 28, 1, 1, 43, -1, 1) op_6947 (v6653[41:0], v6654[27:0], v6947[42:0]); // 7.0
    wire [39:0] v6948; shift_adder #(39, 39, 1, 1, 40, 0, 0) op_6948 (v6655[38:0], v6656[38:0], v6948[39:0]); // 7.0
    wire [36:0] v6949; shift_adder #(36, 35, 1, 1, 37, -1, 0) op_6949 (v6657[35:0], v6658[34:0], v6949[36:0]); // 7.0
    wire [32:0] v6950; shift_adder #(33, 27, 1, 1, 33, 1, 0) op_6950 (v6659[32:0], v6660[26:0], v6950[32:0]); // 7.0
    wire [34:0] v6951; shift_adder #(28, 28, 1, 1, 35, 7, 0) op_6951 (v6661[27:0], v6662[27:0], v6951[34:0]); // 7.0
    wire [36:0] v6952; shift_adder #(34, 34, 1, 1, 37, 2, 0) op_6952 (v6663[33:0], v6664[33:0], v6952[36:0]); // 7.0
    wire [41:0] v6953; shift_adder #(42, 27, 1, 1, 42, 4, 1) op_6953 (v6665[41:0], v6666[26:0], v6953[41:0]); // 7.0
    wire [39:0] v6954; shift_adder #(38, 37, 1, 1, 40, 2, 0) op_6954 (v6667[37:0], v6668[36:0], v6954[39:0]); // 7.0
    wire [36:0] v6955; shift_adder #(36, 35, 1, 1, 37, 0, 0) op_6955 (v6669[35:0], v6670[34:0], v6955[36:0]); // 7.0
    wire [33:0] v6956; shift_adder #(32, 31, 1, 1, 34, -2, 0) op_6956 (v6671[31:0], v6672[30:0], v6956[33:0]); // 7.0
    wire [34:0] v6957; shift_adder #(32, 30, 1, 1, 35, 5, 0) op_6957 (v6673[31:0], v6674[29:0], v6957[34:0]); // 7.0
    wire [34:0] v6958; shift_adder #(27, 27, 1, 1, 35, 8, 1) op_6958 (v6675[26:0], v6127[26:0], v6958[34:0]); // 7.0
    wire [38:0] v6959; shift_adder #(36, 38, 1, 1, 39, -1, 0) op_6959 (v6676[35:0], v6677[37:0], v6959[38:0]); // 7.0
    wire [42:0] v6960; shift_adder #(43, 21, 1, 1, 43, 3, 1) op_6960 (v6678[42:0], v6679[20:0], v6960[42:0]); // 7.0
    wire [31:0] v6961; shift_adder #(31, 30, 1, 1, 32, -1, 0) op_6961 (v6680[30:0], v6681[29:0], v6961[31:0]); // 7.0
    wire [30:0] v6962; shift_adder #(29, 27, 1, 1, 31, -2, 0) op_6962 (v6682[28:0], v6683[26:0], v6962[30:0]); // 7.0
    wire [31:0] v6963; shift_adder #(24, 32, 1, 1, 32, -2, 0) op_6963 (v6684[23:0], v6685[31:0], v6963[31:0]); // 7.0
    wire [32:0] v6964; shift_adder #(33, 29, 1, 1, 33, 0, 0) op_6964 (v6687[32:0], v6625[28:0], v6964[32:0]); // 7.0
    wire [38:0] v6965; shift_adder #(39, 23, 1, 1, 39, 2, 1) op_6965 (v6688[38:0], v6689[22:0], v6965[38:0]); // 7.0
    wire [33:0] v6966; shift_adder #(31, 30, 1, 1, 34, -3, 0) op_6966 (v6690[30:0], v6691[29:0], v6966[33:0]); // 7.0
    wire [34:0] v6967; shift_adder #(33, 34, 1, 1, 35, 1, 0) op_6967 (v6692[32:0], v6693[33:0], v6967[34:0]); // 7.0
    wire [37:0] v6968; shift_adder #(37, 36, 1, 1, 38, 1, 0) op_6968 (v6694[36:0], v6695[35:0], v6968[37:0]); // 7.0
    wire [34:0] v6969; shift_adder #(30, 29, 1, 1, 35, 5, 0) op_6969 (v6696[29:0], v6697[28:0], v6969[34:0]); // 7.0
    wire [35:0] v6970; shift_adder #(35, 33, 1, 1, 36, -1, 0) op_6970 (v6699[34:0], v6700[32:0], v6970[35:0]); // 7.0
    wire [37:0] v6971; shift_adder #(22, 37, 1, 1, 38, 1, 1) op_6971 (v6701[21:0], v6176[36:0], v6971[37:0]); // 7.0
    wire [31:0] v6972; shift_adder #(29, 29, 1, 1, 32, -3, 0) op_6972 (v6702[28:0], v6703[28:0], v6972[31:0]); // 7.0
    wire [41:0] v6973; shift_adder #(39, 36, 1, 1, 42, 5, 0) op_6973 (v6704[38:0], v6705[35:0], v6973[41:0]); // 7.0
    wire [38:0] v6974; shift_adder #(39, 25, 1, 1, 39, 1, 1) op_6974 (v6706[38:0], v6707[24:0], v6974[38:0]); // 7.0
    wire [30:0] v6975; shift_adder #(27, 30, 1, 1, 31, 1, 0) op_6975 (v6708[26:0], v6709[29:0], v6975[30:0]); // 7.0
    wire [34:0] v6976; shift_adder #(33, 31, 1, 1, 35, 3, 0) op_6976 (v6710[32:0], v6711[30:0], v6976[34:0]); // 7.0
    wire [37:0] v6977; shift_adder #(37, 26, 1, 1, 38, -1, 1) op_6977 (v6712[36:0], v6713[25:0], v6977[37:0]); // 7.0
    wire [39:0] v6978; shift_adder #(37, 39, 1, 1, 40, -1, 0) op_6978 (v6714[36:0], v6715[38:0], v6978[39:0]); // 7.0
    wire [32:0] v6979; shift_adder #(31, 32, 1, 1, 33, -2, 0) op_6979 (v6716[30:0], v6717[31:0], v6979[32:0]); // 7.0
    wire [31:0] v6980; shift_adder #(31, 29, 1, 1, 32, 0, 0) op_6980 (v6718[30:0], v6719[28:0], v6980[31:0]); // 7.0
    wire [30:0] v6981; shift_adder #(27, 27, 1, 1, 31, 4, 0) op_6981 (v6720[26:0], v6721[26:0], v6981[30:0]); // 7.0
    wire [34:0] v6982; shift_adder #(31, 34, 1, 1, 35, 1, 0) op_6982 (v6722[30:0], v6723[33:0], v6982[34:0]); // 7.0
    wire [40:0] v6983; shift_adder #(41, 25, 1, 1, 41, 4, 1) op_6983 (v6724[40:0], v6725[24:0], v6983[40:0]); // 7.0
    wire [39:0] v6984; shift_adder #(31, 39, 1, 1, 40, -7, 0) op_6984 (v6606[30:0], v6726[38:0], v6984[39:0]); // 7.0
    wire [35:0] v6985; shift_adder #(35, 34, 1, 1, 36, -1, 0) op_6985 (v6727[34:0], v6728[33:0], v6985[35:0]); // 7.0
    wire [37:0] v6986; shift_adder #(37, 30, 1, 1, 38, 3, 0) op_6986 (v6729[36:0], v6730[29:0], v6986[37:0]); // 7.0
    wire [36:0] v6987; shift_adder #(33, 37, 1, 1, 37, 0, 0) op_6987 (v6731[32:0], v6732[36:0], v6987[36:0]); // 7.0
    wire [37:0] v6988; shift_adder #(27, 37, 1, 1, 38, 1, 1) op_6988 (v6733[26:0], v6238[36:0], v6988[37:0]); // 7.0
    wire [36:0] v6989; shift_adder #(35, 35, 1, 1, 37, 1, 0) op_6989 (v6734[34:0], v6735[34:0], v6989[36:0]); // 7.0
    wire [40:0] v6990; shift_adder #(41, 25, 1, 1, 41, 1, 1) op_6990 (v6736[40:0], v6737[24:0], v6990[40:0]); // 7.0
    wire [36:0] v6991; shift_adder #(36, 34, 1, 1, 37, 2, 0) op_6991 (v6738[35:0], v6739[33:0], v6991[36:0]); // 7.0
    wire [30:0] v6992; shift_adder #(25, 25, 1, 1, 31, -6, 0) op_6992 (v6740[24:0], v6741[24:0], v6992[30:0]); // 7.0
    wire [31:0] v6993; shift_adder #(26, 32, 1, 1, 32, -1, 0) op_6993 (v6742[25:0], v6743[31:0], v6993[31:0]); // 7.0
    wire [32:0] v6994; shift_adder #(28, 33, 1, 1, 33, -1, 0) op_6994 (v6744[27:0], v6745[32:0], v6994[32:0]); // 7.0
    wire [41:0] v6995; shift_adder #(39, 41, 1, 1, 42, -1, 0) op_6995 (v6746[38:0], v6747[40:0], v6995[41:0]); // 7.0
    wire [26:0] v6996; shift_adder #(27, 23, 1, 1, 27, 1, 0) op_6996 (v6748[26:0], v6749[22:0], v6996[26:0]); // 7.0
    wire [33:0] v6997; shift_adder #(32, 31, 1, 1, 34, -2, 0) op_6997 (v6750[31:0], v6751[30:0], v6997[33:0]); // 7.0
    wire [32:0] v6998; shift_adder #(33, 29, 1, 1, 33, 0, 0) op_6998 (v6752[32:0], v6753[28:0], v6998[32:0]); // 7.0
    wire [29:0] v6999; shift_adder #(27, 28, 1, 1, 30, 2, 0) op_6999 (v6754[26:0], v6755[27:0], v6999[29:0]); // 7.0
    wire [37:0] v7000; shift_adder #(31, 38, 1, 1, 38, -3, 0) op_7000 (v6756[30:0], v6757[37:0], v7000[37:0]); // 7.0
    wire [40:0] v7001; shift_adder #(39, 39, 1, 1, 41, 1, 0) op_7001 (v6758[38:0], v6759[38:0], v7001[40:0]); // 7.0
    wire [27:0] v7002; shift_adder #(25, 23, 1, 1, 28, -3, 0) op_7002 (v6760[24:0], v6761[22:0], v7002[27:0]); // 7.0
    wire [36:0] v7003; shift_adder #(37, 35, 1, 1, 37, 1, 0) op_7003 (v6762[36:0], v6763[34:0], v7003[36:0]); // 7.0
    wire [31:0] v7004; shift_adder #(30, 29, 1, 1, 32, -2, 0) op_7004 (v6764[29:0], v6765[28:0], v7004[31:0]); // 7.0
    wire [30:0] v7005; shift_adder #(28, 29, 1, 1, 31, 2, 0) op_7005 (v6766[27:0], v6767[28:0], v7005[30:0]); // 7.0
    wire [35:0] v7006; shift_adder #(32, 35, 1, 1, 36, -1, 0) op_7006 (v6768[31:0], v6769[34:0], v7006[35:0]); // 7.0
    wire [41:0] v7007; shift_adder #(42, 23, 1, 1, 42, 2, 1) op_7007 (v6770[41:0], v6771[22:0], v7007[41:0]); // 7.0
    wire [38:0] v7008; shift_adder #(37, 38, 1, 1, 39, 0, 0) op_7008 (v6772[36:0], v6773[37:0], v7008[38:0]); // 7.0
    wire [33:0] v7009; shift_adder #(34, 32, 1, 1, 34, 0, 0) op_7009 (v6774[33:0], v6775[31:0], v7009[33:0]); // 7.0
    wire [33:0] v7010; shift_adder #(33, 28, 1, 1, 34, -1, 0) op_7010 (v6776[32:0], v6777[27:0], v7010[33:0]); // 7.0
    wire [33:0] v7011; shift_adder #(24, 34, 1, 1, 34, -2, 0) op_7011 (v6778[23:0], v6779[33:0], v7011[33:0]); // 7.0
    wire [39:0] v7012; shift_adder #(35, 40, 1, 1, 40, -3, 0) op_7012 (v6781[34:0], v6782[39:0], v7012[39:0]); // 7.0
    wire [38:0] v7013; shift_adder #(39, 22, 1, 1, 39, 1, 1) op_7013 (v6783[38:0], v6784[21:0], v7013[38:0]); // 7.0
    wire [34:0] v7014; shift_adder #(32, 31, 1, 1, 35, -3, 0) op_7014 (v6785[31:0], v6786[30:0], v7014[34:0]); // 7.0
    wire [29:0] v7015; shift_adder #(30, 26, 1, 1, 30, 1, 0) op_7015 (v6787[29:0], v6788[25:0], v7015[29:0]); // 7.0
    wire [31:0] v7016; shift_adder #(28, 26, 1, 1, 32, 6, 0) op_7016 (v6789[27:0], v6790[25:0], v7016[31:0]); // 7.0
    wire [37:0] v7017; shift_adder #(33, 37, 1, 1, 38, 1, 0) op_7017 (v6791[32:0], v6792[36:0], v7017[37:0]); // 7.0
    wire [38:0] v7018; shift_adder #(39, 26, 1, 1, 39, 0, 1) op_7018 (v6793[38:0], v6794[25:0], v7018[38:0]); // 7.0
    wire [41:0] v7019; shift_adder #(38, 42, 1, 1, 42, -3, 0) op_7019 (v6795[37:0], v6796[41:0], v7019[41:0]); // 7.0
    wire [36:0] v7020; shift_adder #(33, 35, 1, 1, 37, -3, 0) op_7020 (v6797[32:0], v6798[34:0], v7020[36:0]); // 7.0
    wire [32:0] v7021; shift_adder #(33, 29, 1, 1, 33, 1, 0) op_7021 (v6799[32:0], v6800[28:0], v7021[32:0]); // 7.0
    wire [31:0] v7022; shift_adder #(28, 32, 1, 1, 32, -1, 0) op_7022 (v6801[27:0], v6802[31:0], v7022[31:0]); // 7.0
    wire [33:0] v7023; shift_adder #(33, 31, 1, 1, 34, 1, 0) op_7023 (v6700[32:0], v6804[30:0], v7023[33:0]); // 7.0
    wire [37:0] v7024; shift_adder #(35, 36, 1, 1, 38, 2, 0) op_7024 (v6805[34:0], v6806[35:0], v7024[37:0]); // 7.0
    wire [40:0] v7025; shift_adder #(40, 36, 1, 1, 41, 4, 0) op_7025 (v6807[39:0], v6506[35:0], v7025[40:0]); // 7.0
    wire [42:0] v7026; shift_adder #(42, 40, 1, 1, 43, 2, 0) op_7026 (v6808[41:0], v6809[39:0], v7026[42:0]); // 7.0
    wire [30:0] v7027; shift_adder #(31, 23, 1, 1, 31, 0, 0) op_7027 (v6810[30:0], v6811[22:0], v7027[30:0]); // 7.0
    wire [27:0] v7028; shift_adder #(24, 27, 1, 1, 28, 1, 0) op_7028 (v6812[23:0], v6813[26:0], v7028[27:0]); // 7.0
    wire [33:0] v7029; shift_adder #(32, 33, 1, 1, 34, 1, 0) op_7029 (v6814[31:0], v6493[32:0], v7029[33:0]); // 7.0
    wire [39:0] v7030; shift_adder #(32, 40, 1, 1, 40, -4, 0) op_7030 (v6815[31:0], v6816[39:0], v7030[39:0]); // 7.0
    wire [40:0] v7031; shift_adder #(40, 39, 1, 1, 41, 0, 0) op_7031 (v6817[39:0], v6818[38:0], v7031[40:0]); // 7.0
    wire [35:0] v7032; shift_adder #(36, 31, 1, 1, 36, 2, 0) op_7032 (v6819[35:0], v6820[30:0], v7032[35:0]); // 7.0
    wire [30:0] v7033; shift_adder #(29, 26, 1, 1, 31, -2, 0) op_7033 (v6821[28:0], v6822[25:0], v7033[30:0]); // 7.0
    wire [34:0] v7034; shift_adder #(30, 34, 1, 1, 35, -2, 0) op_7034 (v6823[29:0], v6824[33:0], v7034[34:0]); // 7.0
    wire [39:0] v7035; shift_adder #(28, 24, 1, 1, 40, 16, 1) op_7035 (v6825[27:0], v6410[23:0], v7035[39:0]); // 7.0
    wire [40:0] v7036; shift_adder #(41, 24, 1, 1, 41, 2, 1) op_7036 (v6826[40:0], v6827[23:0], v7036[40:0]); // 7.0
    wire [42:0] v7037; shift_adder #(42, 36, 1, 1, 43, 6, 0) op_7037 (v6828[41:0], v6829[35:0], v7037[42:0]); // 7.0
    wire [35:0] v7038; shift_adder #(36, 32, 1, 1, 36, 0, 0) op_7038 (v6830[35:0], v6831[31:0], v7038[35:0]); // 7.0
    wire [32:0] v7039; shift_adder #(33, 29, 1, 1, 33, 2, 0) op_7039 (v6832[32:0], v6833[28:0], v7039[32:0]); // 7.0
    wire [29:0] v7040; shift_adder #(22, 28, 1, 1, 30, 2, 0) op_7040 (v6834[21:0], v6835[27:0], v7040[29:0]); // 7.0
    wire [34:0] v7041; shift_adder #(33, 35, 1, 1, 35, 0, 0) op_7041 (v6837[32:0], v6838[34:0], v7041[34:0]); // 7.0
    wire [39:0] v7042; shift_adder #(33, 40, 1, 1, 40, -4, 0) op_7042 (v6839[32:0], v6840[39:0], v7042[39:0]); // 7.0
    wire [35:0] v7043; shift_adder #(33, 32, 1, 1, 36, -3, 0) op_7043 (v6841[32:0], v6842[31:0], v7043[35:0]); // 7.0
    wire [26:0] v7044; shift_adder #(27, 20, 1, 1, 27, 0, 0) op_7044 (v6843[26:0], v6844[19:0], v7044[26:0]); // 7.0
    wire [27:0] v7045; shift_adder #(24, 26, 1, 1, 28, 2, 0) op_7045 (v6845[23:0], v6846[25:0], v7045[27:0]); // 7.0
    wire [33:0] v7046; shift_adder #(32, 33, 1, 1, 34, 1, 0) op_7046 (v6848[31:0], v6849[32:0], v7046[33:0]); // 7.0
    wire [42:0] v7047; shift_adder #(36, 42, 1, 1, 43, -6, 0) op_7047 (v6850[35:0], v6851[41:0], v7047[42:0]); // 7.0
    wire [36:0] v7048; shift_adder #(35, 32, 1, 1, 37, -1, 0) op_7048 (v6852[34:0], v6853[31:0], v7048[36:0]); // 7.0
    wire [28:0] v7049; shift_adder #(29, 25, 1, 1, 29, 0, 0) op_7049 (v6854[28:0], v6855[24:0], v7049[28:0]); // 7.0
    wire [35:0] v7050; shift_adder #(34, 31, 1, 1, 36, 5, 0) op_7050 (v6856[33:0], v6857[30:0], v7050[35:0]); // 7.0
    wire [38:0] v7051; shift_adder #(27, 31, 1, 1, 39, 8, 1) op_7051 (v6858[26:0], v6475[30:0], v7051[38:0]); // 7.0
    wire [39:0] v7052; shift_adder #(34, 39, 1, 1, 40, -3, 0) op_7052 (v6859[33:0], v6860[38:0], v7052[39:0]); // 7.0
    wire [39:0] v7053; shift_adder #(38, 38, 1, 1, 40, 1, 0) op_7053 (v6861[37:0], v6862[37:0], v7053[39:0]); // 7.0
    wire [39:0] v7054; shift_adder #(39, 31, 1, 1, 40, 6, 0) op_7054 (v6863[38:0], v6864[30:0], v7054[39:0]); // 7.0
    wire [34:0] v7055; shift_adder #(35, 27, 1, 1, 35, 3, 0) op_7055 (v6865[34:0], v6866[26:0], v7055[34:0]); // 7.0
    wire [33:0] v7056; shift_adder #(30, 34, 1, 1, 34, 0, 0) op_7056 (v6867[29:0], v6868[33:0], v7056[33:0]); // 8.0
    wire [39:0] v7057; shift_adder #(39, 40, 1, 1, 40, 0, 0) op_7057 (v6870[38:0], v6871[39:0], v7057[39:0]); // 8.0
    wire [39:0] v7058; shift_adder #(38, 33, 1, 1, 40, -2, 1) op_7058 (v6872[37:0], v6873[32:0], v7058[39:0]); // 8.0
    wire [36:0] v7059; shift_adder #(32, 36, 1, 1, 37, 1, 1) op_7059 (v6874[31:0], v6506[35:0], v7059[36:0]); // 8.0
    wire [38:0] v7060; shift_adder #(36, 38, 1, 1, 39, -2, 0) op_7060 (v6876[35:0], v6877[37:0], v7060[38:0]); // 8.0
    wire [40:0] v7061; shift_adder #(41, 32, 1, 1, 41, 3, 1) op_7061 (v6878[40:0], v6879[31:0], v7061[40:0]); // 8.0
    wire [39:0] v7062; shift_adder #(34, 37, 1, 1, 40, 3, 1) op_7062 (v6880[33:0], v6519[36:0], v7062[39:0]); // 8.0
    wire [42:0] v7063; shift_adder #(41, 32, 1, 1, 43, -2, 1) op_7063 (v6882[40:0], v6883[31:0], v7063[42:0]); // 8.0
    wire [43:0] v7064; shift_adder #(36, 44, 1, 1, 44, -6, 0) op_7064 (v6884[35:0], v6885[43:0], v7064[43:0]); // 8.0
    wire [39:0] v7065; shift_adder #(29, 40, 1, 1, 40, -3, 0) op_7065 (v6886[28:0], v6887[39:0], v7065[39:0]); // 8.0
    wire [39:0] v7066; shift_adder #(39, 34, 1, 1, 40, -1, 1) op_7066 (v6888[38:0], v6889[33:0], v7066[39:0]); // 8.0
    wire [39:0] v7067; shift_adder #(40, 36, 1, 1, 40, 1, 0) op_7067 (v6890[39:0], v6891[35:0], v7067[39:0]); // 8.0
    wire [38:0] v7068; shift_adder #(34, 36, 1, 1, 39, 3, 0) op_7068 (v6892[33:0], v6893[35:0], v7068[38:0]); // 8.0
    wire [41:0] v7069; shift_adder #(39, 42, 1, 1, 42, -2, 0) op_7069 (v6894[38:0], v6895[41:0], v7069[41:0]); // 8.0
    wire [36:0] v7070; shift_adder #(37, 30, 1, 1, 37, 0, 0) op_7070 (v6896[36:0], v6897[29:0], v7070[36:0]); // 8.0
    wire [43:0] v7071; shift_adder #(37, 22, 1, 1, 44, 22, 1) op_7071 (v6898[36:0], v6555[21:0], v7071[43:0]); // 8.0
    wire [40:0] v7072; shift_adder #(38, 33, 1, 1, 41, -3, 1) op_7072 (v6900[37:0], v6901[32:0], v7072[40:0]); // 8.0
    wire [41:0] v7073; shift_adder #(37, 42, 1, 1, 42, -2, 0) op_7073 (v6902[36:0], v6903[41:0], v7073[41:0]); // 8.0
    wire [35:0] v7074; shift_adder #(28, 35, 1, 1, 36, 1, 0) op_7074 (v6904[27:0], v6905[34:0], v7074[35:0]); // 8.0
    wire [42:0] v7075; shift_adder #(41, 41, 1, 1, 43, 2, 0) op_7075 (v6906[40:0], v6907[40:0], v7075[42:0]); // 8.0
    wire [36:0] v7076; shift_adder #(37, 31, 1, 1, 37, 0, 0) op_7076 (v6908[36:0], v6909[30:0], v7076[36:0]); // 8.0
    wire [39:0] v7077; shift_adder #(32, 40, 1, 1, 40, -1, 0) op_7077 (v6910[31:0], v6911[39:0], v7077[39:0]); // 8.0
    wire [39:0] v7078; shift_adder #(39, 31, 1, 1, 40, -1, 1) op_7078 (v6912[38:0], v6913[30:0], v7078[39:0]); // 8.0
    wire [36:0] v7079; shift_adder #(34, 32, 1, 1, 37, -3, 0) op_7079 (v6914[33:0], v6915[31:0], v7079[36:0]); // 8.0
    wire [32:0] v7080; shift_adder #(30, 28, 1, 1, 33, 5, 1) op_7080 (v6916[29:0], v6592[27:0], v7080[32:0]); // 8.0
    wire [40:0] v7081; shift_adder #(40, 39, 1, 1, 41, 1, 0) op_7081 (v6918[39:0], v6919[38:0], v7081[40:0]); // 8.0
    wire [41:0] v7082; shift_adder #(39, 42, 1, 1, 42, -2, 0) op_7082 (v6920[38:0], v6921[41:0], v7082[41:0]); // 8.0
    wire [36:0] v7083; shift_adder #(31, 30, 1, 1, 37, 7, 0) op_7083 (v6922[30:0], v6923[29:0], v7083[36:0]); // 8.0
    wire [41:0] v7084; shift_adder #(37, 42, 1, 1, 42, -2, 0) op_7084 (v6924[36:0], v6925[41:0], v7084[41:0]); // 8.0
    wire [42:0] v7085; shift_adder #(37, 35, 1, 1, 43, -6, 0) op_7085 (v6926[36:0], v6927[34:0], v7085[42:0]); // 8.0
    wire [40:0] v7086; shift_adder #(32, 36, 1, 1, 41, 5, 1) op_7086 (v6928[31:0], v6616[35:0], v7086[40:0]); // 8.0
    wire [41:0] v7087; shift_adder #(40, 42, 1, 1, 42, 0, 0) op_7087 (v6929[39:0], v6930[41:0], v7087[41:0]); // 8.0
    wire [37:0] v7088; shift_adder #(36, 32, 1, 1, 38, -2, 0) op_7088 (v6931[35:0], v6932[31:0], v7088[37:0]); // 8.0
    wire [35:0] v7089; shift_adder #(31, 36, 1, 1, 36, -2, 1) op_7089 (v6933[30:0], v6627[35:0], v7089[35:0]); // 8.0
    wire [39:0] v7090; shift_adder #(38, 38, 1, 1, 40, 2, 0) op_7090 (v6935[37:0], v6936[37:0], v7090[39:0]); // 8.0
    wire [41:0] v7091; shift_adder #(41, 41, 1, 1, 42, 0, 0) op_7091 (v6937[40:0], v6938[40:0], v7091[41:0]); // 8.0
    wire [37:0] v7092; shift_adder #(32, 38, 1, 1, 38, 0, 0) op_7092 (v6939[31:0], v6940[37:0], v7092[37:0]); // 8.0
    wire [41:0] v7093; shift_adder #(42, 27, 1, 1, 42, 3, 1) op_7093 (v6941[41:0], v6942[26:0], v7093[41:0]); // 8.0
    wire [35:0] v7094; shift_adder #(36, 33, 1, 1, 36, 0, 0) op_7094 (v6943[35:0], v6944[32:0], v7094[35:0]); // 8.0
    wire [37:0] v7095; shift_adder #(32, 37, 1, 1, 38, 1, 0) op_7095 (v6945[31:0], v6946[36:0], v7095[37:0]); // 8.0
    wire [44:0] v7096; shift_adder #(43, 40, 1, 1, 45, 4, 0) op_7096 (v6947[42:0], v6948[39:0], v7096[44:0]); // 8.0
    wire [37:0] v7097; shift_adder #(37, 33, 1, 1, 38, -1, 0) op_7097 (v6949[36:0], v6950[32:0], v7097[37:0]); // 8.0
    wire [40:0] v7098; shift_adder #(35, 37, 1, 1, 41, 4, 0) op_7098 (v6951[34:0], v6952[36:0], v7098[40:0]); // 8.0
    wire [42:0] v7099; shift_adder #(42, 40, 1, 1, 43, 2, 0) op_7099 (v6953[41:0], v6954[39:0], v7099[42:0]); // 8.0
    wire [37:0] v7100; shift_adder #(37, 34, 1, 1, 38, -1, 0) op_7100 (v6955[36:0], v6956[33:0], v7100[37:0]); // 8.0
    wire [36:0] v7101; shift_adder #(35, 35, 1, 1, 37, 1, 0) op_7101 (v6957[34:0], v6958[34:0], v7101[36:0]); // 8.0
    wire [42:0] v7102; shift_adder #(39, 43, 1, 1, 43, -3, 0) op_7102 (v6959[38:0], v6960[42:0], v7102[42:0]); // 8.0
    wire [36:0] v7103; shift_adder #(32, 31, 1, 1, 37, -5, 0) op_7103 (v6961[31:0], v6962[30:0], v7103[36:0]); // 8.0
    wire [39:0] v7104; shift_adder #(32, 38, 1, 1, 40, 2, 1) op_7104 (v6963[31:0], v6686[37:0], v7104[39:0]); // 8.0
    wire [40:0] v7105; shift_adder #(39, 34, 1, 1, 41, -2, 1) op_7105 (v6965[38:0], v6966[33:0], v7105[40:0]); // 8.0
    wire [37:0] v7106; shift_adder #(35, 38, 1, 1, 38, -1, 0) op_7106 (v6967[34:0], v6968[37:0], v7106[37:0]); // 8.0
    wire [39:0] v7107; shift_adder #(35, 29, 1, 1, 40, 11, 1) op_7107 (v6969[34:0], v6698[28:0], v7107[39:0]); // 8.0
    wire [38:0] v7108; shift_adder #(38, 32, 1, 1, 39, -1, 1) op_7108 (v6971[37:0], v6972[31:0], v7108[38:0]); // 8.0
    wire [41:0] v7109; shift_adder #(42, 39, 1, 1, 42, 2, 0) op_7109 (v6973[41:0], v6974[38:0], v7109[41:0]); // 8.0
    wire [37:0] v7110; shift_adder #(31, 35, 1, 1, 38, 3, 0) op_7110 (v6975[30:0], v6976[34:0], v7110[37:0]); // 8.0
    wire [39:0] v7111; shift_adder #(38, 40, 1, 1, 40, -1, 0) op_7111 (v6977[37:0], v6978[39:0], v7111[39:0]); // 8.0
    wire [36:0] v7112; shift_adder #(33, 32, 1, 1, 37, -4, 0) op_7112 (v6979[32:0], v6980[31:0], v7112[36:0]); // 8.0
    wire [37:0] v7113; shift_adder #(31, 35, 1, 1, 38, 3, 0) op_7113 (v6981[30:0], v6982[34:0], v7113[37:0]); // 8.0
    wire [41:0] v7114; shift_adder #(41, 40, 1, 1, 42, 1, 0) op_7114 (v6983[40:0], v6984[39:0], v7114[41:0]); // 8.0
    wire [40:0] v7115; shift_adder #(36, 38, 1, 1, 41, -4, 0) op_7115 (v6985[35:0], v6986[37:0], v7115[40:0]); // 8.0
    wire [38:0] v7116; shift_adder #(37, 38, 1, 1, 39, 1, 0) op_7116 (v6987[36:0], v6988[37:0], v7116[38:0]); // 8.0
    wire [41:0] v7117; shift_adder #(37, 41, 1, 1, 42, -4, 0) op_7117 (v6989[36:0], v6990[40:0], v7117[41:0]); // 8.0
    wire [36:0] v7118; shift_adder #(37, 31, 1, 1, 37, 0, 0) op_7118 (v6991[36:0], v6992[30:0], v7118[36:0]); // 8.0
    wire [39:0] v7119; shift_adder #(32, 33, 1, 1, 40, 7, 0) op_7119 (v6993[31:0], v6994[32:0], v7119[39:0]); // 8.0
    wire [41:0] v7120; shift_adder #(42, 27, 1, 1, 42, 1, 1) op_7120 (v6995[41:0], v6996[26:0], v7120[41:0]); // 8.0
    wire [36:0] v7121; shift_adder #(34, 33, 1, 1, 37, -3, 0) op_7121 (v6997[33:0], v6998[32:0], v7121[36:0]); // 8.0
    wire [37:0] v7122; shift_adder #(30, 38, 1, 1, 38, 0, 0) op_7122 (v6999[29:0], v7000[37:0], v7122[37:0]); // 8.0
    wire [40:0] v7123; shift_adder #(41, 28, 1, 1, 41, 1, 1) op_7123 (v7001[40:0], v7002[27:0], v7123[40:0]); // 8.0
    wire [37:0] v7124; shift_adder #(37, 32, 1, 1, 38, 1, 0) op_7124 (v7003[36:0], v7004[31:0], v7124[37:0]); // 8.0
    wire [36:0] v7125; shift_adder #(31, 36, 1, 1, 37, 1, 0) op_7125 (v7005[30:0], v7006[35:0], v7125[36:0]); // 8.0
    wire [42:0] v7126; shift_adder #(42, 39, 1, 1, 43, 4, 0) op_7126 (v7007[41:0], v7008[38:0], v7126[42:0]); // 8.0
    wire [36:0] v7127; shift_adder #(34, 34, 1, 1, 37, -2, 0) op_7127 (v7009[33:0], v7010[33:0], v7127[36:0]); // 8.0
    wire [40:0] v7128; shift_adder #(34, 33, 1, 1, 41, 8, 1) op_7128 (v7011[33:0], v6780[32:0], v7128[40:0]); // 8.0
    wire [41:0] v7129; shift_adder #(40, 39, 1, 1, 42, 3, 0) op_7129 (v7012[39:0], v7013[38:0], v7129[41:0]); // 8.0
    wire [35:0] v7130; shift_adder #(35, 30, 1, 1, 36, -1, 0) op_7130 (v7014[34:0], v7015[29:0], v7130[35:0]); // 8.0
    wire [38:0] v7131; shift_adder #(32, 38, 1, 1, 39, 1, 0) op_7131 (v7016[31:0], v7017[37:0], v7131[38:0]); // 8.0
    wire [42:0] v7132; shift_adder #(39, 42, 1, 1, 43, -2, 0) op_7132 (v7018[38:0], v7019[41:0], v7132[42:0]); // 8.0
    wire [38:0] v7133; shift_adder #(37, 33, 1, 1, 39, -2, 0) op_7133 (v7020[36:0], v7021[32:0], v7133[38:0]); // 8.0
    wire [38:0] v7134; shift_adder #(32, 30, 1, 1, 39, 9, 1) op_7134 (v7022[31:0], v6803[29:0], v7134[38:0]); // 8.0
    wire [40:0] v7135; shift_adder #(38, 41, 1, 1, 41, -1, 0) op_7135 (v7024[37:0], v7025[40:0], v7135[40:0]); // 8.0
    wire [42:0] v7136; shift_adder #(43, 31, 1, 1, 43, 3, 1) op_7136 (v7026[42:0], v7027[30:0], v7136[42:0]); // 8.0
    wire [35:0] v7137; shift_adder #(28, 34, 1, 1, 36, 2, 0) op_7137 (v7028[27:0], v7029[33:0], v7137[35:0]); // 8.0
    wire [40:0] v7138; shift_adder #(40, 41, 1, 1, 41, 0, 0) op_7138 (v7030[39:0], v7031[40:0], v7138[40:0]); // 8.0
    wire [38:0] v7139; shift_adder #(36, 31, 1, 1, 39, -3, 0) op_7139 (v7032[35:0], v7033[30:0], v7139[38:0]); // 8.0
    wire [39:0] v7140; shift_adder #(35, 40, 1, 1, 40, -3, 0) op_7140 (v7034[34:0], v7035[39:0], v7140[39:0]); // 8.0
    wire [43:0] v7141; shift_adder #(41, 43, 1, 1, 44, -2, 0) op_7141 (v7036[40:0], v7037[42:0], v7141[43:0]); // 8.0
    wire [39:0] v7142; shift_adder #(36, 33, 1, 1, 40, -4, 0) op_7142 (v7038[35:0], v7039[32:0], v7142[39:0]); // 8.0
    wire [40:0] v7143; shift_adder #(30, 34, 1, 1, 41, 7, 1) op_7143 (v7040[29:0], v6836[33:0], v7143[40:0]); // 8.0
    wire [39:0] v7144; shift_adder #(35, 40, 1, 1, 40, 0, 0) op_7144 (v7041[34:0], v7042[39:0], v7144[39:0]); // 8.0
    wire [35:0] v7145; shift_adder #(36, 27, 1, 1, 36, 1, 0) op_7145 (v7043[35:0], v7044[26:0], v7145[35:0]); // 8.0
    wire [39:0] v7146; shift_adder #(28, 34, 1, 1, 40, 6, 1) op_7146 (v7045[27:0], v6847[33:0], v7146[39:0]); // 8.0
    wire [42:0] v7147; shift_adder #(34, 43, 1, 1, 43, -4, 0) op_7147 (v7046[33:0], v7047[42:0], v7147[42:0]); // 8.0
    wire [39:0] v7148; shift_adder #(37, 29, 1, 1, 40, -3, 0) op_7148 (v7048[36:0], v7049[28:0], v7148[39:0]); // 8.0
    wire [38:0] v7149; shift_adder #(36, 39, 1, 1, 39, -1, 0) op_7149 (v7050[35:0], v7051[38:0], v7149[38:0]); // 8.0
    wire [40:0] v7150; shift_adder #(40, 40, 1, 1, 41, 1, 0) op_7150 (v7052[39:0], v7053[39:0], v7150[40:0]); // 8.0
    wire [40:0] v7151; shift_adder #(40, 35, 1, 1, 41, -1, 0) op_7151 (v7054[39:0], v7055[34:0], v7151[40:0]); // 8.0
    wire [35:0] v7152; shift_adder #(34, 35, 1, 1, 36, 0, 1) op_7152 (v7056[33:0], v6869[34:0], v7152[35:0]); // 9.0
    wire [40:0] v7153; shift_adder #(40, 40, 1, 1, 41, 0, 0) op_7153 (v7057[39:0], v7058[39:0], v7153[40:0]); // 9.0
    wire [37:0] v7154; shift_adder #(37, 33, 1, 1, 38, 5, 1) op_7154 (v7059[36:0], v6875[32:0], v7154[37:0]); // 9.0
    wire [41:0] v7155; shift_adder #(39, 41, 1, 1, 42, -2, 0) op_7155 (v7060[38:0], v7061[40:0], v7155[41:0]); // 9.0
    wire [39:0] v7156; shift_adder #(40, 34, 1, 1, 40, 4, 1) op_7156 (v7062[39:0], v6881[33:0], v7156[39:0]); // 9.0
    wire [44:0] v7157; shift_adder #(43, 44, 1, 1, 45, -1, 0) op_7157 (v7063[42:0], v7064[43:0], v7157[44:0]); // 9.0
    wire [41:0] v7158; shift_adder #(40, 40, 1, 1, 42, 2, 0) op_7158 (v7065[39:0], v7066[39:0], v7158[41:0]); // 9.0
    wire [41:0] v7159; shift_adder #(39, 42, 1, 1, 42, 0, 0) op_7159 (v7068[38:0], v7069[41:0], v7159[41:0]); // 9.0
    wire [44:0] v7160; shift_adder #(44, 38, 1, 1, 45, 6, 1) op_7160 (v7071[43:0], v6899[37:0], v7160[44:0]); // 9.0
    wire [42:0] v7161; shift_adder #(41, 42, 1, 1, 43, -1, 0) op_7161 (v7072[40:0], v7073[41:0], v7161[42:0]); // 9.0
    wire [42:0] v7162; shift_adder #(36, 43, 1, 1, 43, -3, 0) op_7162 (v7074[35:0], v7075[42:0], v7162[42:0]); // 9.0
    wire [41:0] v7163; shift_adder #(40, 40, 1, 1, 42, 1, 0) op_7163 (v7077[39:0], v7078[39:0], v7163[41:0]); // 9.0
    wire [35:0] v7164; shift_adder #(33, 31, 1, 1, 36, -3, 1) op_7164 (v7080[32:0], v6917[30:0], v7164[35:0]); // 9.0
    wire [42:0] v7165; shift_adder #(41, 42, 1, 1, 43, 0, 0) op_7165 (v7081[40:0], v7082[41:0], v7165[42:0]); // 9.0
    wire [41:0] v7166; shift_adder #(37, 42, 1, 1, 42, 0, 0) op_7166 (v7083[36:0], v7084[41:0], v7166[41:0]); // 9.0
    wire [42:0] v7167; shift_adder #(41, 42, 1, 1, 43, 0, 0) op_7167 (v7086[40:0], v7087[41:0], v7167[42:0]); // 9.0
    wire [36:0] v7168; shift_adder #(36, 35, 1, 1, 37, -1, 1) op_7168 (v7089[35:0], v6934[34:0], v7168[36:0]); // 9.0
    wire [42:0] v7169; shift_adder #(40, 42, 1, 1, 43, 0, 0) op_7169 (v7090[39:0], v7091[41:0], v7169[42:0]); // 9.0
    wire [41:0] v7170; shift_adder #(38, 42, 1, 1, 42, -2, 0) op_7170 (v7092[37:0], v7093[41:0], v7170[41:0]); // 9.0
    wire [44:0] v7171; shift_adder #(38, 45, 1, 1, 45, -4, 0) op_7171 (v7095[37:0], v7096[44:0], v7171[44:0]); // 9.0
    wire [43:0] v7172; shift_adder #(41, 43, 1, 1, 44, 1, 0) op_7172 (v7098[40:0], v7099[42:0], v7172[43:0]); // 9.0
    wire [42:0] v7173; shift_adder #(37, 43, 1, 1, 43, -4, 0) op_7173 (v7101[36:0], v7102[42:0], v7173[42:0]); // 9.0
    wire [39:0] v7174; shift_adder #(40, 33, 1, 1, 40, 3, 1) op_7174 (v7104[39:0], v6964[32:0], v7174[39:0]); // 9.0
    wire [41:0] v7175; shift_adder #(41, 38, 1, 1, 42, 3, 0) op_7175 (v7105[40:0], v7106[37:0], v7175[41:0]); // 9.0
    wire [40:0] v7176; shift_adder #(40, 36, 1, 1, 41, 3, 1) op_7176 (v7107[39:0], v6970[35:0], v7176[40:0]); // 9.0
    wire [42:0] v7177; shift_adder #(39, 42, 1, 1, 43, -3, 0) op_7177 (v7108[38:0], v7109[41:0], v7177[42:0]); // 9.0
    wire [40:0] v7178; shift_adder #(38, 40, 1, 1, 41, 0, 0) op_7178 (v7110[37:0], v7111[39:0], v7178[40:0]); // 9.0
    wire [41:0] v7179; shift_adder #(38, 42, 1, 1, 42, 0, 0) op_7179 (v7113[37:0], v7114[41:0], v7179[41:0]); // 9.0
    wire [41:0] v7180; shift_adder #(39, 42, 1, 1, 42, -1, 0) op_7180 (v7116[38:0], v7117[41:0], v7180[41:0]); // 9.0
    wire [41:0] v7181; shift_adder #(40, 42, 1, 1, 42, 0, 0) op_7181 (v7119[39:0], v7120[41:0], v7181[41:0]); // 9.0
    wire [40:0] v7182; shift_adder #(38, 41, 1, 1, 41, -1, 0) op_7182 (v7122[37:0], v7123[40:0], v7182[40:0]); // 9.0
    wire [42:0] v7183; shift_adder #(37, 43, 1, 1, 43, -3, 0) op_7183 (v7125[36:0], v7126[42:0], v7183[42:0]); // 9.0
    wire [42:0] v7184; shift_adder #(41, 42, 1, 1, 43, 0, 0) op_7184 (v7128[40:0], v7129[41:0], v7184[42:0]); // 9.0
    wire [42:0] v7185; shift_adder #(39, 43, 1, 1, 43, -1, 0) op_7185 (v7131[38:0], v7132[42:0], v7185[42:0]); // 9.0
    wire [38:0] v7186; shift_adder #(39, 34, 1, 1, 39, 4, 1) op_7186 (v7134[38:0], v7023[33:0], v7186[38:0]); // 9.0
    wire [42:0] v7187; shift_adder #(41, 43, 1, 1, 43, 0, 0) op_7187 (v7135[40:0], v7136[42:0], v7187[42:0]); // 9.0
    wire [40:0] v7188; shift_adder #(36, 41, 1, 1, 41, -1, 0) op_7188 (v7137[35:0], v7138[40:0], v7188[40:0]); // 9.0
    wire [44:0] v7189; shift_adder #(40, 44, 1, 1, 45, -3, 0) op_7189 (v7140[39:0], v7141[43:0], v7189[44:0]); // 9.0
    wire [42:0] v7190; shift_adder #(41, 40, 1, 1, 43, 2, 0) op_7190 (v7143[40:0], v7144[39:0], v7190[42:0]); // 9.0
    wire [43:0] v7191; shift_adder #(40, 43, 1, 1, 44, -2, 0) op_7191 (v7146[39:0], v7147[42:0], v7191[43:0]); // 9.0
    wire [41:0] v7192; shift_adder #(39, 41, 1, 1, 42, 1, 0) op_7192 (v7149[38:0], v7150[40:0], v7192[41:0]); // 9.0
    wire [41:0] v7193; shift_adder #(36, 41, 1, 1, 42, -4, 0) op_7193 (v7152[35:0], v7153[40:0], v7193[41:0]); // 10.0
    wire [42:0] v7194; shift_adder #(38, 42, 1, 1, 43, -3, 0) op_7194 (v7154[37:0], v7155[41:0], v7194[42:0]); // 10.0
    wire [45:0] v7195; shift_adder #(40, 45, 1, 1, 46, -3, 0) op_7195 (v7156[39:0], v7157[44:0], v7195[45:0]); // 10.0
    wire [43:0] v7196; shift_adder #(42, 40, 1, 1, 44, 3, 1) op_7196 (v7158[41:0], v7067[39:0], v7196[43:0]); // 10.0
    wire [42:0] v7197; shift_adder #(42, 37, 1, 1, 43, 4, 1) op_7197 (v7159[41:0], v7070[36:0], v7197[42:0]); // 10.0
    wire [46:0] v7198; shift_adder #(45, 43, 1, 1, 47, 3, 0) op_7198 (v7160[44:0], v7161[42:0], v7198[46:0]); // 10.0
    wire [43:0] v7199; shift_adder #(43, 37, 1, 1, 44, 5, 1) op_7199 (v7162[42:0], v7076[36:0], v7199[43:0]); // 10.0
    wire [41:0] v7200; shift_adder #(42, 37, 1, 1, 42, 4, 1) op_7200 (v7163[41:0], v7079[36:0], v7200[41:0]); // 10.0
    wire [42:0] v7201; shift_adder #(36, 43, 1, 1, 43, -2, 0) op_7201 (v7164[35:0], v7165[42:0], v7201[42:0]); // 10.0
    wire [44:0] v7202; shift_adder #(42, 43, 1, 1, 45, -2, 1) op_7202 (v7166[41:0], v7085[42:0], v7202[44:0]); // 10.0
    wire [42:0] v7203; shift_adder #(43, 38, 1, 1, 43, 2, 1) op_7203 (v7167[42:0], v7088[37:0], v7203[42:0]); // 10.0
    wire [42:0] v7204; shift_adder #(37, 43, 1, 1, 43, -1, 0) op_7204 (v7168[36:0], v7169[42:0], v7204[42:0]); // 10.0
    wire [42:0] v7205; shift_adder #(42, 36, 1, 1, 43, 5, 1) op_7205 (v7170[41:0], v7094[35:0], v7205[42:0]); // 10.0
    wire [45:0] v7206; shift_adder #(45, 38, 1, 1, 46, 6, 1) op_7206 (v7171[44:0], v7097[37:0], v7206[45:0]); // 10.0
    wire [44:0] v7207; shift_adder #(44, 38, 1, 1, 45, 5, 1) op_7207 (v7172[43:0], v7100[37:0], v7207[44:0]); // 10.0
    wire [43:0] v7208; shift_adder #(43, 37, 1, 1, 44, 3, 1) op_7208 (v7173[42:0], v7103[36:0], v7208[43:0]); // 10.0
    wire [42:0] v7209; shift_adder #(40, 42, 1, 1, 43, -1, 0) op_7209 (v7174[39:0], v7175[41:0], v7209[42:0]); // 10.0
    wire [43:0] v7210; shift_adder #(41, 43, 1, 1, 44, -1, 0) op_7210 (v7176[40:0], v7177[42:0], v7210[43:0]); // 10.0
    wire [40:0] v7211; shift_adder #(41, 37, 1, 1, 41, 1, 1) op_7211 (v7178[40:0], v7112[36:0], v7211[40:0]); // 10.0
    wire [42:0] v7212; shift_adder #(42, 41, 1, 1, 43, 1, 1) op_7212 (v7179[41:0], v7115[40:0], v7212[42:0]); // 10.0
    wire [42:0] v7213; shift_adder #(42, 37, 1, 1, 43, 4, 1) op_7213 (v7180[41:0], v7118[36:0], v7213[42:0]); // 10.0
    wire [42:0] v7214; shift_adder #(42, 37, 1, 1, 43, 4, 1) op_7214 (v7181[41:0], v7121[36:0], v7214[42:0]); // 10.0
    wire [41:0] v7215; shift_adder #(41, 38, 1, 1, 42, 3, 1) op_7215 (v7182[40:0], v7124[37:0], v7215[41:0]); // 10.0
    wire [43:0] v7216; shift_adder #(43, 37, 1, 1, 44, 5, 1) op_7216 (v7183[42:0], v7127[36:0], v7216[43:0]); // 10.0
    wire [42:0] v7217; shift_adder #(43, 36, 1, 1, 43, 3, 1) op_7217 (v7184[42:0], v7130[35:0], v7217[42:0]); // 10.0
    wire [43:0] v7218; shift_adder #(43, 39, 1, 1, 44, 3, 1) op_7218 (v7185[42:0], v7133[38:0], v7218[43:0]); // 10.0
    wire [43:0] v7219; shift_adder #(39, 43, 1, 1, 44, -2, 0) op_7219 (v7186[38:0], v7187[42:0], v7219[43:0]); // 10.0
    wire [41:0] v7220; shift_adder #(41, 39, 1, 1, 42, 1, 1) op_7220 (v7188[40:0], v7139[38:0], v7220[41:0]); // 10.0
    wire [44:0] v7221; shift_adder #(45, 40, 1, 1, 45, 2, 1) op_7221 (v7189[44:0], v7142[39:0], v7221[44:0]); // 10.0
    wire [42:0] v7222; shift_adder #(43, 36, 1, 1, 43, 2, 1) op_7222 (v7190[42:0], v7145[35:0], v7222[42:0]); // 10.0
    wire [43:0] v7223; shift_adder #(44, 40, 1, 1, 44, 1, 1) op_7223 (v7191[43:0], v7148[39:0], v7223[43:0]); // 10.0
    wire [43:0] v7224; shift_adder #(42, 41, 1, 1, 44, -1, 1) op_7224 (v7192[41:0], v7151[40:0], v7224[43:0]); // 10.0

    // verilator lint_on UNUSEDSIGNAL

    assign out[41:0] = v7193[41:0];
    assign out[84:42] = v7194[42:0];
    assign out[130:85] = v7195[45:0];
    assign out[174:131] = v7196[43:0];
    assign out[217:175] = v7197[42:0];
    assign out[264:218] = v7198[46:0];
    assign out[308:265] = v7199[43:0];
    assign out[350:309] = v7200[41:0];
    assign out[393:351] = v7201[42:0];
    assign out[438:394] = v7202[44:0];
    assign out[481:439] = v7203[42:0];
    assign out[524:482] = v7204[42:0];
    assign out[567:525] = v7205[42:0];
    assign out[613:568] = v7206[45:0];
    assign out[658:614] = v7207[44:0];
    assign out[702:659] = v7208[43:0];
    assign out[745:703] = v7209[42:0];
    assign out[789:746] = v7210[43:0];
    assign out[830:790] = v7211[40:0];
    assign out[873:831] = v7212[42:0];
    assign out[916:874] = v7213[42:0];
    assign out[959:917] = v7214[42:0];
    assign out[1001:960] = v7215[41:0];
    assign out[1045:1002] = v7216[43:0];
    assign out[1088:1046] = v7217[42:0];
    assign out[1132:1089] = v7218[43:0];
    assign out[1176:1133] = v7219[43:0];
    assign out[1218:1177] = v7220[41:0];
    assign out[1263:1219] = v7221[44:0];
    assign out[1306:1264] = v7222[42:0];
    assign out[1350:1307] = v7223[43:0];
    assign out[1394:1351] = v7224[43:0];

    endmodule
